VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_counter
  CLASS BLOCK ;
  FOREIGN wrapped_counter ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.300 4.000 12.500 ;
    END
  END active
  PIN chip_pin_output_bit[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 246.000 14.770 250.000 ;
    END
  END chip_pin_output_bit[0]
  PIN chip_pin_output_bit[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.810 246.000 42.370 250.000 ;
    END
  END chip_pin_output_bit[1]
  PIN chip_pin_output_bit[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.410 246.000 69.970 250.000 ;
    END
  END chip_pin_output_bit[2]
  PIN chip_pin_output_bit[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 246.000 97.570 250.000 ;
    END
  END chip_pin_output_bit[3]
  PIN chip_pin_output_bit[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.610 246.000 125.170 250.000 ;
    END
  END chip_pin_output_bit[4]
  PIN chip_pin_output_bit[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.210 246.000 152.770 250.000 ;
    END
  END chip_pin_output_bit[5]
  PIN chip_pin_output_bit[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 246.000 180.370 250.000 ;
    END
  END chip_pin_output_bit[6]
  PIN chip_pin_output_bit[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.410 246.000 207.970 250.000 ;
    END
  END chip_pin_output_bit[7]
  PIN clk_blip
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.010 246.000 235.570 250.000 ;
    END
  END clk_blip
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.420 4.000 18.620 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.620 4.000 79.820 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.740 4.000 85.940 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.860 4.000 92.060 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.980 4.000 98.180 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.100 4.000 104.300 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.220 4.000 110.420 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.340 4.000 116.540 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.460 4.000 122.660 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.580 4.000 128.780 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.700 4.000 134.900 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.540 4.000 24.740 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.820 4.000 141.020 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.940 4.000 147.140 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.060 4.000 153.260 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.180 4.000 159.380 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.300 4.000 165.500 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.420 4.000 171.620 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.540 4.000 177.740 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.660 4.000 183.860 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.780 4.000 189.980 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.900 4.000 196.100 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.660 4.000 30.860 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.020 4.000 202.220 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.140 4.000 208.340 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.260 4.000 214.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.380 4.000 220.580 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.500 4.000 226.700 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.620 4.000 232.820 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.740 4.000 238.940 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.860 4.000 245.060 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.780 4.000 36.980 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.900 4.000 43.100 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.020 4.000 49.220 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.140 4.000 55.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.260 4.000 61.460 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.380 4.000 67.580 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.500 4.000 73.700 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.990 0.000 126.550 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.190 0.000 158.750 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.410 0.000 161.970 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.630 0.000 165.190 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 0.000 168.410 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.070 0.000 171.630 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.290 0.000 174.850 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.510 0.000 178.070 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.730 0.000 181.290 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.950 0.000 184.510 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.170 0.000 187.730 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.210 0.000 129.770 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.390 0.000 190.950 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.610 0.000 194.170 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.830 0.000 197.390 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.050 0.000 200.610 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 0.000 203.830 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.490 0.000 207.050 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.710 0.000 210.270 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.930 0.000 213.490 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.150 0.000 216.710 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.370 0.000 219.930 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 0.000 132.990 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.590 0.000 223.150 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.810 0.000 226.370 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.030 0.000 229.590 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.250 0.000 232.810 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.470 0.000 236.030 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.690 0.000 239.250 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.910 0.000 242.470 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.130 0.000 245.690 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.650 0.000 136.210 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.870 0.000 139.430 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.090 0.000 142.650 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.310 0.000 145.870 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.530 0.000 149.090 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.750 0.000 152.310 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.970 0.000 155.530 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.630 0.000 4.190 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.830 0.000 36.390 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.050 0.000 39.610 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.270 0.000 42.830 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.490 0.000 46.050 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.710 0.000 49.270 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.930 0.000 52.490 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.150 0.000 55.710 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.370 0.000 58.930 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 0.000 62.150 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.810 0.000 65.370 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.850 0.000 7.410 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.030 0.000 68.590 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.250 0.000 71.810 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.470 0.000 75.030 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.690 0.000 78.250 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.910 0.000 81.470 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.130 0.000 84.690 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.350 0.000 87.910 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.570 0.000 91.130 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.790 0.000 94.350 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 0.000 97.570 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.070 0.000 10.630 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.230 0.000 100.790 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.450 0.000 104.010 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.670 0.000 107.230 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.890 0.000 110.450 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.110 0.000 113.670 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.330 0.000 116.890 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.550 0.000 120.110 4.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.770 0.000 123.330 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.290 0.000 13.850 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.510 0.000 17.070 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.730 0.000 20.290 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.950 0.000 23.510 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 0.000 26.730 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.390 0.000 29.950 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.610 0.000 33.170 4.000 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 236.880 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.180 4.000 6.380 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 244.260 236.725 ;
      LAYER met1 ;
        RECT 3.750 6.840 245.570 236.880 ;
      LAYER met2 ;
        RECT 3.780 245.720 13.930 246.570 ;
        RECT 15.050 245.720 41.530 246.570 ;
        RECT 42.650 245.720 69.130 246.570 ;
        RECT 70.250 245.720 96.730 246.570 ;
        RECT 97.850 245.720 124.330 246.570 ;
        RECT 125.450 245.720 151.930 246.570 ;
        RECT 153.050 245.720 179.530 246.570 ;
        RECT 180.650 245.720 207.130 246.570 ;
        RECT 208.250 245.720 234.730 246.570 ;
        RECT 235.850 245.720 245.540 246.570 ;
        RECT 3.780 4.280 245.540 245.720 ;
        RECT 4.470 4.000 6.570 4.280 ;
        RECT 7.690 4.000 9.790 4.280 ;
        RECT 10.910 4.000 13.010 4.280 ;
        RECT 14.130 4.000 16.230 4.280 ;
        RECT 17.350 4.000 19.450 4.280 ;
        RECT 20.570 4.000 22.670 4.280 ;
        RECT 23.790 4.000 25.890 4.280 ;
        RECT 27.010 4.000 29.110 4.280 ;
        RECT 30.230 4.000 32.330 4.280 ;
        RECT 33.450 4.000 35.550 4.280 ;
        RECT 36.670 4.000 38.770 4.280 ;
        RECT 39.890 4.000 41.990 4.280 ;
        RECT 43.110 4.000 45.210 4.280 ;
        RECT 46.330 4.000 48.430 4.280 ;
        RECT 49.550 4.000 51.650 4.280 ;
        RECT 52.770 4.000 54.870 4.280 ;
        RECT 55.990 4.000 58.090 4.280 ;
        RECT 59.210 4.000 61.310 4.280 ;
        RECT 62.430 4.000 64.530 4.280 ;
        RECT 65.650 4.000 67.750 4.280 ;
        RECT 68.870 4.000 70.970 4.280 ;
        RECT 72.090 4.000 74.190 4.280 ;
        RECT 75.310 4.000 77.410 4.280 ;
        RECT 78.530 4.000 80.630 4.280 ;
        RECT 81.750 4.000 83.850 4.280 ;
        RECT 84.970 4.000 87.070 4.280 ;
        RECT 88.190 4.000 90.290 4.280 ;
        RECT 91.410 4.000 93.510 4.280 ;
        RECT 94.630 4.000 96.730 4.280 ;
        RECT 97.850 4.000 99.950 4.280 ;
        RECT 101.070 4.000 103.170 4.280 ;
        RECT 104.290 4.000 106.390 4.280 ;
        RECT 107.510 4.000 109.610 4.280 ;
        RECT 110.730 4.000 112.830 4.280 ;
        RECT 113.950 4.000 116.050 4.280 ;
        RECT 117.170 4.000 119.270 4.280 ;
        RECT 120.390 4.000 122.490 4.280 ;
        RECT 123.610 4.000 125.710 4.280 ;
        RECT 126.830 4.000 128.930 4.280 ;
        RECT 130.050 4.000 132.150 4.280 ;
        RECT 133.270 4.000 135.370 4.280 ;
        RECT 136.490 4.000 138.590 4.280 ;
        RECT 139.710 4.000 141.810 4.280 ;
        RECT 142.930 4.000 145.030 4.280 ;
        RECT 146.150 4.000 148.250 4.280 ;
        RECT 149.370 4.000 151.470 4.280 ;
        RECT 152.590 4.000 154.690 4.280 ;
        RECT 155.810 4.000 157.910 4.280 ;
        RECT 159.030 4.000 161.130 4.280 ;
        RECT 162.250 4.000 164.350 4.280 ;
        RECT 165.470 4.000 167.570 4.280 ;
        RECT 168.690 4.000 170.790 4.280 ;
        RECT 171.910 4.000 174.010 4.280 ;
        RECT 175.130 4.000 177.230 4.280 ;
        RECT 178.350 4.000 180.450 4.280 ;
        RECT 181.570 4.000 183.670 4.280 ;
        RECT 184.790 4.000 186.890 4.280 ;
        RECT 188.010 4.000 190.110 4.280 ;
        RECT 191.230 4.000 193.330 4.280 ;
        RECT 194.450 4.000 196.550 4.280 ;
        RECT 197.670 4.000 199.770 4.280 ;
        RECT 200.890 4.000 202.990 4.280 ;
        RECT 204.110 4.000 206.210 4.280 ;
        RECT 207.330 4.000 209.430 4.280 ;
        RECT 210.550 4.000 212.650 4.280 ;
        RECT 213.770 4.000 215.870 4.280 ;
        RECT 216.990 4.000 219.090 4.280 ;
        RECT 220.210 4.000 222.310 4.280 ;
        RECT 223.430 4.000 225.530 4.280 ;
        RECT 226.650 4.000 228.750 4.280 ;
        RECT 229.870 4.000 231.970 4.280 ;
        RECT 233.090 4.000 235.190 4.280 ;
        RECT 236.310 4.000 238.410 4.280 ;
        RECT 239.530 4.000 241.630 4.280 ;
        RECT 242.750 4.000 244.850 4.280 ;
      LAYER met3 ;
        RECT 4.000 233.220 176.230 236.805 ;
        RECT 4.400 231.220 176.230 233.220 ;
        RECT 4.000 227.100 176.230 231.220 ;
        RECT 4.400 225.100 176.230 227.100 ;
        RECT 4.000 220.980 176.230 225.100 ;
        RECT 4.400 218.980 176.230 220.980 ;
        RECT 4.000 214.860 176.230 218.980 ;
        RECT 4.400 212.860 176.230 214.860 ;
        RECT 4.000 208.740 176.230 212.860 ;
        RECT 4.400 206.740 176.230 208.740 ;
        RECT 4.000 202.620 176.230 206.740 ;
        RECT 4.400 200.620 176.230 202.620 ;
        RECT 4.000 196.500 176.230 200.620 ;
        RECT 4.400 194.500 176.230 196.500 ;
        RECT 4.000 190.380 176.230 194.500 ;
        RECT 4.400 188.380 176.230 190.380 ;
        RECT 4.000 184.260 176.230 188.380 ;
        RECT 4.400 182.260 176.230 184.260 ;
        RECT 4.000 178.140 176.230 182.260 ;
        RECT 4.400 176.140 176.230 178.140 ;
        RECT 4.000 172.020 176.230 176.140 ;
        RECT 4.400 170.020 176.230 172.020 ;
        RECT 4.000 165.900 176.230 170.020 ;
        RECT 4.400 163.900 176.230 165.900 ;
        RECT 4.000 159.780 176.230 163.900 ;
        RECT 4.400 157.780 176.230 159.780 ;
        RECT 4.000 153.660 176.230 157.780 ;
        RECT 4.400 151.660 176.230 153.660 ;
        RECT 4.000 147.540 176.230 151.660 ;
        RECT 4.400 145.540 176.230 147.540 ;
        RECT 4.000 141.420 176.230 145.540 ;
        RECT 4.400 139.420 176.230 141.420 ;
        RECT 4.000 135.300 176.230 139.420 ;
        RECT 4.400 133.300 176.230 135.300 ;
        RECT 4.000 129.180 176.230 133.300 ;
        RECT 4.400 127.180 176.230 129.180 ;
        RECT 4.000 123.060 176.230 127.180 ;
        RECT 4.400 121.060 176.230 123.060 ;
        RECT 4.000 116.940 176.230 121.060 ;
        RECT 4.400 114.940 176.230 116.940 ;
        RECT 4.000 110.820 176.230 114.940 ;
        RECT 4.400 108.820 176.230 110.820 ;
        RECT 4.000 104.700 176.230 108.820 ;
        RECT 4.400 102.700 176.230 104.700 ;
        RECT 4.000 98.580 176.230 102.700 ;
        RECT 4.400 96.580 176.230 98.580 ;
        RECT 4.000 92.460 176.230 96.580 ;
        RECT 4.400 90.460 176.230 92.460 ;
        RECT 4.000 86.340 176.230 90.460 ;
        RECT 4.400 84.340 176.230 86.340 ;
        RECT 4.000 80.220 176.230 84.340 ;
        RECT 4.400 78.220 176.230 80.220 ;
        RECT 4.000 74.100 176.230 78.220 ;
        RECT 4.400 72.100 176.230 74.100 ;
        RECT 4.000 67.980 176.230 72.100 ;
        RECT 4.400 65.980 176.230 67.980 ;
        RECT 4.000 61.860 176.230 65.980 ;
        RECT 4.400 59.860 176.230 61.860 ;
        RECT 4.000 55.740 176.230 59.860 ;
        RECT 4.400 53.740 176.230 55.740 ;
        RECT 4.000 49.620 176.230 53.740 ;
        RECT 4.400 47.620 176.230 49.620 ;
        RECT 4.000 43.500 176.230 47.620 ;
        RECT 4.400 41.500 176.230 43.500 ;
        RECT 4.000 37.380 176.230 41.500 ;
        RECT 4.400 35.380 176.230 37.380 ;
        RECT 4.000 31.260 176.230 35.380 ;
        RECT 4.400 29.260 176.230 31.260 ;
        RECT 4.000 25.140 176.230 29.260 ;
        RECT 4.400 23.140 176.230 25.140 ;
        RECT 4.000 19.020 176.230 23.140 ;
        RECT 4.400 17.020 176.230 19.020 ;
        RECT 4.000 12.900 176.230 17.020 ;
        RECT 4.400 10.900 176.230 12.900 ;
        RECT 4.000 10.715 176.230 10.900 ;
  END
END wrapped_counter
END LIBRARY

