module wrapper_squared
(
  output wire [37:0] io_out,
  output wire [37:0] io_oeb,
  inout wire vccd1,
  inout wire vcca1,
  inout wire vssa1,
  inout wire vssd1,
  inout wire [10:0] analog_io,
  input wire wb_clk_i,
  input wire [37:0] io_in,
  input wire active
);

endmodule
