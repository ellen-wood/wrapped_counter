magic
tech sky130B
magscale 1 2
timestamp 1672306177
<< obsli1 >>
rect 1104 2159 48852 47345
<< obsm1 >>
rect 750 1504 49114 47376
<< metal2 >>
rect 1738 49200 1850 50000
rect 5050 49200 5162 50000
rect 8362 49200 8474 50000
rect 11674 49200 11786 50000
rect 14986 49200 15098 50000
rect 18298 49200 18410 50000
rect 21610 49200 21722 50000
rect 24922 49200 25034 50000
rect 28234 49200 28346 50000
rect 31546 49200 31658 50000
rect 34858 49200 34970 50000
rect 38170 49200 38282 50000
rect 41482 49200 41594 50000
rect 44794 49200 44906 50000
rect 48106 49200 48218 50000
rect 726 0 838 800
rect 1370 0 1482 800
rect 2014 0 2126 800
rect 2658 0 2770 800
rect 3302 0 3414 800
rect 3946 0 4058 800
rect 4590 0 4702 800
rect 5234 0 5346 800
rect 5878 0 5990 800
rect 6522 0 6634 800
rect 7166 0 7278 800
rect 7810 0 7922 800
rect 8454 0 8566 800
rect 9098 0 9210 800
rect 9742 0 9854 800
rect 10386 0 10498 800
rect 11030 0 11142 800
rect 11674 0 11786 800
rect 12318 0 12430 800
rect 12962 0 13074 800
rect 13606 0 13718 800
rect 14250 0 14362 800
rect 14894 0 15006 800
rect 15538 0 15650 800
rect 16182 0 16294 800
rect 16826 0 16938 800
rect 17470 0 17582 800
rect 18114 0 18226 800
rect 18758 0 18870 800
rect 19402 0 19514 800
rect 20046 0 20158 800
rect 20690 0 20802 800
rect 21334 0 21446 800
rect 21978 0 22090 800
rect 22622 0 22734 800
rect 23266 0 23378 800
rect 23910 0 24022 800
rect 24554 0 24666 800
rect 25198 0 25310 800
rect 25842 0 25954 800
rect 26486 0 26598 800
rect 27130 0 27242 800
rect 27774 0 27886 800
rect 28418 0 28530 800
rect 29062 0 29174 800
rect 29706 0 29818 800
rect 30350 0 30462 800
rect 30994 0 31106 800
rect 31638 0 31750 800
rect 32282 0 32394 800
rect 32926 0 33038 800
rect 33570 0 33682 800
rect 34214 0 34326 800
rect 34858 0 34970 800
rect 35502 0 35614 800
rect 36146 0 36258 800
rect 36790 0 36902 800
rect 37434 0 37546 800
rect 38078 0 38190 800
rect 38722 0 38834 800
rect 39366 0 39478 800
rect 40010 0 40122 800
rect 40654 0 40766 800
rect 41298 0 41410 800
rect 41942 0 42054 800
rect 42586 0 42698 800
rect 43230 0 43342 800
rect 43874 0 43986 800
rect 44518 0 44630 800
rect 45162 0 45274 800
rect 45806 0 45918 800
rect 46450 0 46562 800
rect 47094 0 47206 800
rect 47738 0 47850 800
rect 48382 0 48494 800
rect 49026 0 49138 800
<< obsm2 >>
rect 756 49144 1682 49314
rect 1906 49144 4994 49314
rect 5218 49144 8306 49314
rect 8530 49144 11618 49314
rect 11842 49144 14930 49314
rect 15154 49144 18242 49314
rect 18466 49144 21554 49314
rect 21778 49144 24866 49314
rect 25090 49144 28178 49314
rect 28402 49144 31490 49314
rect 31714 49144 34802 49314
rect 35026 49144 38114 49314
rect 38338 49144 41426 49314
rect 41650 49144 44738 49314
rect 44962 49144 48050 49314
rect 48274 49144 49108 49314
rect 756 856 49108 49144
rect 894 800 1314 856
rect 1538 800 1958 856
rect 2182 800 2602 856
rect 2826 800 3246 856
rect 3470 800 3890 856
rect 4114 800 4534 856
rect 4758 800 5178 856
rect 5402 800 5822 856
rect 6046 800 6466 856
rect 6690 800 7110 856
rect 7334 800 7754 856
rect 7978 800 8398 856
rect 8622 800 9042 856
rect 9266 800 9686 856
rect 9910 800 10330 856
rect 10554 800 10974 856
rect 11198 800 11618 856
rect 11842 800 12262 856
rect 12486 800 12906 856
rect 13130 800 13550 856
rect 13774 800 14194 856
rect 14418 800 14838 856
rect 15062 800 15482 856
rect 15706 800 16126 856
rect 16350 800 16770 856
rect 16994 800 17414 856
rect 17638 800 18058 856
rect 18282 800 18702 856
rect 18926 800 19346 856
rect 19570 800 19990 856
rect 20214 800 20634 856
rect 20858 800 21278 856
rect 21502 800 21922 856
rect 22146 800 22566 856
rect 22790 800 23210 856
rect 23434 800 23854 856
rect 24078 800 24498 856
rect 24722 800 25142 856
rect 25366 800 25786 856
rect 26010 800 26430 856
rect 26654 800 27074 856
rect 27298 800 27718 856
rect 27942 800 28362 856
rect 28586 800 29006 856
rect 29230 800 29650 856
rect 29874 800 30294 856
rect 30518 800 30938 856
rect 31162 800 31582 856
rect 31806 800 32226 856
rect 32450 800 32870 856
rect 33094 800 33514 856
rect 33738 800 34158 856
rect 34382 800 34802 856
rect 35026 800 35446 856
rect 35670 800 36090 856
rect 36314 800 36734 856
rect 36958 800 37378 856
rect 37602 800 38022 856
rect 38246 800 38666 856
rect 38890 800 39310 856
rect 39534 800 39954 856
rect 40178 800 40598 856
rect 40822 800 41242 856
rect 41466 800 41886 856
rect 42110 800 42530 856
rect 42754 800 43174 856
rect 43398 800 43818 856
rect 44042 800 44462 856
rect 44686 800 45106 856
rect 45330 800 45750 856
rect 45974 800 46394 856
rect 46618 800 47038 856
rect 47262 800 47682 856
rect 47906 800 48326 856
rect 48550 800 48970 856
<< metal3 >>
rect 0 47276 800 47516
rect 0 45916 800 46156
rect 0 44556 800 44796
rect 0 43196 800 43436
rect 0 41836 800 42076
rect 0 40476 800 40716
rect 0 39116 800 39356
rect 0 37756 800 37996
rect 0 36396 800 36636
rect 0 35036 800 35276
rect 0 33676 800 33916
rect 0 32316 800 32556
rect 0 30956 800 31196
rect 0 29596 800 29836
rect 0 28236 800 28476
rect 0 26876 800 27116
rect 0 25516 800 25756
rect 0 24156 800 24396
rect 0 22796 800 23036
rect 0 21436 800 21676
rect 0 20076 800 20316
rect 0 18716 800 18956
rect 0 17356 800 17596
rect 0 15996 800 16236
rect 0 14636 800 14876
rect 0 13276 800 13516
rect 0 11916 800 12156
rect 0 10556 800 10796
rect 0 9196 800 9436
rect 0 7836 800 8076
rect 0 6476 800 6716
rect 0 5116 800 5356
rect 0 3756 800 3996
rect 0 2396 800 2636
<< obsm3 >>
rect 3049 2143 35246 47361
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
<< labels >>
rlabel metal2 s 1738 49200 1850 50000 6 active
port 1 nsew signal input
rlabel metal2 s 21610 49200 21722 50000 6 chip_pin_output_bit[0]
port 2 nsew signal input
rlabel metal2 s 24922 49200 25034 50000 6 chip_pin_output_bit[1]
port 3 nsew signal input
rlabel metal2 s 28234 49200 28346 50000 6 chip_pin_output_bit[2]
port 4 nsew signal input
rlabel metal2 s 31546 49200 31658 50000 6 chip_pin_output_bit[3]
port 5 nsew signal input
rlabel metal2 s 34858 49200 34970 50000 6 chip_pin_output_bit[4]
port 6 nsew signal input
rlabel metal2 s 38170 49200 38282 50000 6 chip_pin_output_bit[5]
port 7 nsew signal input
rlabel metal2 s 41482 49200 41594 50000 6 chip_pin_output_bit[6]
port 8 nsew signal input
rlabel metal2 s 44794 49200 44906 50000 6 chip_pin_output_bit[7]
port 9 nsew signal input
rlabel metal2 s 48106 49200 48218 50000 6 clk_blip
port 10 nsew signal input
rlabel metal3 s 0 3756 800 3996 6 io_in[0]
port 11 nsew signal input
rlabel metal2 s 11674 49200 11786 50000 6 io_in[10]
port 12 nsew signal input
rlabel metal2 s 14986 49200 15098 50000 6 io_in[11]
port 13 nsew signal input
rlabel metal2 s 18298 49200 18410 50000 6 io_in[12]
port 14 nsew signal input
rlabel metal3 s 0 14636 800 14876 6 io_in[13]
port 15 nsew signal input
rlabel metal3 s 0 15996 800 16236 6 io_in[14]
port 16 nsew signal input
rlabel metal3 s 0 17356 800 17596 6 io_in[15]
port 17 nsew signal input
rlabel metal3 s 0 18716 800 18956 6 io_in[16]
port 18 nsew signal input
rlabel metal3 s 0 20076 800 20316 6 io_in[17]
port 19 nsew signal input
rlabel metal3 s 0 21436 800 21676 6 io_in[18]
port 20 nsew signal input
rlabel metal3 s 0 22796 800 23036 6 io_in[19]
port 21 nsew signal input
rlabel metal3 s 0 5116 800 5356 6 io_in[1]
port 22 nsew signal input
rlabel metal3 s 0 24156 800 24396 6 io_in[20]
port 23 nsew signal input
rlabel metal3 s 0 25516 800 25756 6 io_in[21]
port 24 nsew signal input
rlabel metal3 s 0 26876 800 27116 6 io_in[22]
port 25 nsew signal input
rlabel metal3 s 0 28236 800 28476 6 io_in[23]
port 26 nsew signal input
rlabel metal3 s 0 29596 800 29836 6 io_in[24]
port 27 nsew signal input
rlabel metal3 s 0 30956 800 31196 6 io_in[25]
port 28 nsew signal input
rlabel metal3 s 0 32316 800 32556 6 io_in[26]
port 29 nsew signal input
rlabel metal3 s 0 33676 800 33916 6 io_in[27]
port 30 nsew signal input
rlabel metal3 s 0 35036 800 35276 6 io_in[28]
port 31 nsew signal input
rlabel metal3 s 0 36396 800 36636 6 io_in[29]
port 32 nsew signal input
rlabel metal3 s 0 6476 800 6716 6 io_in[2]
port 33 nsew signal input
rlabel metal3 s 0 37756 800 37996 6 io_in[30]
port 34 nsew signal input
rlabel metal3 s 0 39116 800 39356 6 io_in[31]
port 35 nsew signal input
rlabel metal3 s 0 40476 800 40716 6 io_in[32]
port 36 nsew signal input
rlabel metal3 s 0 41836 800 42076 6 io_in[33]
port 37 nsew signal input
rlabel metal3 s 0 43196 800 43436 6 io_in[34]
port 38 nsew signal input
rlabel metal3 s 0 44556 800 44796 6 io_in[35]
port 39 nsew signal input
rlabel metal3 s 0 45916 800 46156 6 io_in[36]
port 40 nsew signal input
rlabel metal3 s 0 47276 800 47516 6 io_in[37]
port 41 nsew signal input
rlabel metal3 s 0 7836 800 8076 6 io_in[3]
port 42 nsew signal input
rlabel metal3 s 0 9196 800 9436 6 io_in[4]
port 43 nsew signal input
rlabel metal3 s 0 10556 800 10796 6 io_in[5]
port 44 nsew signal input
rlabel metal3 s 0 11916 800 12156 6 io_in[6]
port 45 nsew signal input
rlabel metal3 s 0 13276 800 13516 6 io_in[7]
port 46 nsew signal input
rlabel metal2 s 5050 49200 5162 50000 6 io_in[8]
port 47 nsew signal input
rlabel metal2 s 8362 49200 8474 50000 6 io_in[9]
port 48 nsew signal input
rlabel metal2 s 25198 0 25310 800 6 io_oeb[0]
port 49 nsew signal output
rlabel metal2 s 31638 0 31750 800 6 io_oeb[10]
port 50 nsew signal output
rlabel metal2 s 32282 0 32394 800 6 io_oeb[11]
port 51 nsew signal output
rlabel metal2 s 32926 0 33038 800 6 io_oeb[12]
port 52 nsew signal output
rlabel metal2 s 33570 0 33682 800 6 io_oeb[13]
port 53 nsew signal output
rlabel metal2 s 34214 0 34326 800 6 io_oeb[14]
port 54 nsew signal output
rlabel metal2 s 34858 0 34970 800 6 io_oeb[15]
port 55 nsew signal output
rlabel metal2 s 35502 0 35614 800 6 io_oeb[16]
port 56 nsew signal output
rlabel metal2 s 36146 0 36258 800 6 io_oeb[17]
port 57 nsew signal output
rlabel metal2 s 36790 0 36902 800 6 io_oeb[18]
port 58 nsew signal output
rlabel metal2 s 37434 0 37546 800 6 io_oeb[19]
port 59 nsew signal output
rlabel metal2 s 25842 0 25954 800 6 io_oeb[1]
port 60 nsew signal output
rlabel metal2 s 38078 0 38190 800 6 io_oeb[20]
port 61 nsew signal output
rlabel metal2 s 38722 0 38834 800 6 io_oeb[21]
port 62 nsew signal output
rlabel metal2 s 39366 0 39478 800 6 io_oeb[22]
port 63 nsew signal output
rlabel metal2 s 40010 0 40122 800 6 io_oeb[23]
port 64 nsew signal output
rlabel metal2 s 40654 0 40766 800 6 io_oeb[24]
port 65 nsew signal output
rlabel metal2 s 41298 0 41410 800 6 io_oeb[25]
port 66 nsew signal output
rlabel metal2 s 41942 0 42054 800 6 io_oeb[26]
port 67 nsew signal output
rlabel metal2 s 42586 0 42698 800 6 io_oeb[27]
port 68 nsew signal output
rlabel metal2 s 43230 0 43342 800 6 io_oeb[28]
port 69 nsew signal output
rlabel metal2 s 43874 0 43986 800 6 io_oeb[29]
port 70 nsew signal output
rlabel metal2 s 26486 0 26598 800 6 io_oeb[2]
port 71 nsew signal output
rlabel metal2 s 44518 0 44630 800 6 io_oeb[30]
port 72 nsew signal output
rlabel metal2 s 45162 0 45274 800 6 io_oeb[31]
port 73 nsew signal output
rlabel metal2 s 45806 0 45918 800 6 io_oeb[32]
port 74 nsew signal output
rlabel metal2 s 46450 0 46562 800 6 io_oeb[33]
port 75 nsew signal output
rlabel metal2 s 47094 0 47206 800 6 io_oeb[34]
port 76 nsew signal output
rlabel metal2 s 47738 0 47850 800 6 io_oeb[35]
port 77 nsew signal output
rlabel metal2 s 48382 0 48494 800 6 io_oeb[36]
port 78 nsew signal output
rlabel metal2 s 49026 0 49138 800 6 io_oeb[37]
port 79 nsew signal output
rlabel metal2 s 27130 0 27242 800 6 io_oeb[3]
port 80 nsew signal output
rlabel metal2 s 27774 0 27886 800 6 io_oeb[4]
port 81 nsew signal output
rlabel metal2 s 28418 0 28530 800 6 io_oeb[5]
port 82 nsew signal output
rlabel metal2 s 29062 0 29174 800 6 io_oeb[6]
port 83 nsew signal output
rlabel metal2 s 29706 0 29818 800 6 io_oeb[7]
port 84 nsew signal output
rlabel metal2 s 30350 0 30462 800 6 io_oeb[8]
port 85 nsew signal output
rlabel metal2 s 30994 0 31106 800 6 io_oeb[9]
port 86 nsew signal output
rlabel metal2 s 726 0 838 800 6 io_out[0]
port 87 nsew signal output
rlabel metal2 s 7166 0 7278 800 6 io_out[10]
port 88 nsew signal output
rlabel metal2 s 7810 0 7922 800 6 io_out[11]
port 89 nsew signal output
rlabel metal2 s 8454 0 8566 800 6 io_out[12]
port 90 nsew signal output
rlabel metal2 s 9098 0 9210 800 6 io_out[13]
port 91 nsew signal output
rlabel metal2 s 9742 0 9854 800 6 io_out[14]
port 92 nsew signal output
rlabel metal2 s 10386 0 10498 800 6 io_out[15]
port 93 nsew signal output
rlabel metal2 s 11030 0 11142 800 6 io_out[16]
port 94 nsew signal output
rlabel metal2 s 11674 0 11786 800 6 io_out[17]
port 95 nsew signal output
rlabel metal2 s 12318 0 12430 800 6 io_out[18]
port 96 nsew signal output
rlabel metal2 s 12962 0 13074 800 6 io_out[19]
port 97 nsew signal output
rlabel metal2 s 1370 0 1482 800 6 io_out[1]
port 98 nsew signal output
rlabel metal2 s 13606 0 13718 800 6 io_out[20]
port 99 nsew signal output
rlabel metal2 s 14250 0 14362 800 6 io_out[21]
port 100 nsew signal output
rlabel metal2 s 14894 0 15006 800 6 io_out[22]
port 101 nsew signal output
rlabel metal2 s 15538 0 15650 800 6 io_out[23]
port 102 nsew signal output
rlabel metal2 s 16182 0 16294 800 6 io_out[24]
port 103 nsew signal output
rlabel metal2 s 16826 0 16938 800 6 io_out[25]
port 104 nsew signal output
rlabel metal2 s 17470 0 17582 800 6 io_out[26]
port 105 nsew signal output
rlabel metal2 s 18114 0 18226 800 6 io_out[27]
port 106 nsew signal output
rlabel metal2 s 18758 0 18870 800 6 io_out[28]
port 107 nsew signal output
rlabel metal2 s 19402 0 19514 800 6 io_out[29]
port 108 nsew signal output
rlabel metal2 s 2014 0 2126 800 6 io_out[2]
port 109 nsew signal output
rlabel metal2 s 20046 0 20158 800 6 io_out[30]
port 110 nsew signal output
rlabel metal2 s 20690 0 20802 800 6 io_out[31]
port 111 nsew signal output
rlabel metal2 s 21334 0 21446 800 6 io_out[32]
port 112 nsew signal output
rlabel metal2 s 21978 0 22090 800 6 io_out[33]
port 113 nsew signal output
rlabel metal2 s 22622 0 22734 800 6 io_out[34]
port 114 nsew signal output
rlabel metal2 s 23266 0 23378 800 6 io_out[35]
port 115 nsew signal output
rlabel metal2 s 23910 0 24022 800 6 io_out[36]
port 116 nsew signal output
rlabel metal2 s 24554 0 24666 800 6 io_out[37]
port 117 nsew signal output
rlabel metal2 s 2658 0 2770 800 6 io_out[3]
port 118 nsew signal output
rlabel metal2 s 3302 0 3414 800 6 io_out[4]
port 119 nsew signal output
rlabel metal2 s 3946 0 4058 800 6 io_out[5]
port 120 nsew signal output
rlabel metal2 s 4590 0 4702 800 6 io_out[6]
port 121 nsew signal output
rlabel metal2 s 5234 0 5346 800 6 io_out[7]
port 122 nsew signal output
rlabel metal2 s 5878 0 5990 800 6 io_out[8]
port 123 nsew signal output
rlabel metal2 s 6522 0 6634 800 6 io_out[9]
port 124 nsew signal output
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 125 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 125 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 126 nsew ground bidirectional
rlabel metal3 s 0 2396 800 2636 6 wb_clk_i
port 127 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1110856
string GDS_FILE /openlane/designs/wrapped_counter/runs/RUN_2022.12.29_09.28.34/results/signoff/wrapped_counter.magic.gds
string GDS_START 149560
<< end >>

