magic
tech sky130B
magscale 1 2
timestamp 1672306175
<< viali >>
rect 2053 47141 2087 47175
rect 35173 47141 35207 47175
rect 1869 47005 1903 47039
rect 5273 47005 5307 47039
rect 21833 47005 21867 47039
rect 25053 47005 25087 47039
rect 28365 47005 28399 47039
rect 32137 47005 32171 47039
rect 34989 47005 35023 47039
rect 38301 47005 38335 47039
rect 45477 47005 45511 47039
rect 47685 47005 47719 47039
rect 5641 46937 5675 46971
rect 42901 46937 42935 46971
rect 47961 46937 47995 46971
rect 22017 46869 22051 46903
rect 25237 46869 25271 46903
rect 28549 46869 28583 46903
rect 32321 46869 32355 46903
rect 38485 46869 38519 46903
rect 42993 46869 43027 46903
rect 45569 46869 45603 46903
rect 10333 8925 10367 8959
rect 12541 8925 12575 8959
rect 10425 8789 10459 8823
rect 12633 8789 12667 8823
rect 7665 8449 7699 8483
rect 8401 8449 8435 8483
rect 9045 8449 9079 8483
rect 9689 8449 9723 8483
rect 47869 8449 47903 8483
rect 1869 8313 1903 8347
rect 7757 8313 7791 8347
rect 8493 8313 8527 8347
rect 9137 8313 9171 8347
rect 9781 8313 9815 8347
rect 47961 8313 47995 8347
rect 10333 8041 10367 8075
rect 2605 7905 2639 7939
rect 1869 7837 1903 7871
rect 6101 7837 6135 7871
rect 7021 7837 7055 7871
rect 8217 7837 8251 7871
rect 9413 7837 9447 7871
rect 10517 7837 10551 7871
rect 10977 7837 11011 7871
rect 47133 7837 47167 7871
rect 47593 7837 47627 7871
rect 8401 7769 8435 7803
rect 10057 7769 10091 7803
rect 6193 7701 6227 7735
rect 7113 7701 7147 7735
rect 9505 7701 9539 7735
rect 11069 7701 11103 7735
rect 47685 7701 47719 7735
rect 1961 7361 1995 7395
rect 4997 7361 5031 7395
rect 5641 7361 5675 7395
rect 6745 7361 6779 7395
rect 7205 7361 7239 7395
rect 7941 7361 7975 7395
rect 10701 7361 10735 7395
rect 11529 7361 11563 7395
rect 47593 7361 47627 7395
rect 8217 7293 8251 7327
rect 47685 7293 47719 7327
rect 6561 7225 6595 7259
rect 11621 7225 11655 7259
rect 47041 7225 47075 7259
rect 2053 7157 2087 7191
rect 3341 7157 3375 7191
rect 5089 7157 5123 7191
rect 5733 7157 5767 7191
rect 7297 7157 7331 7191
rect 9689 7157 9723 7191
rect 10793 7157 10827 7191
rect 46397 7157 46431 7191
rect 5438 6953 5472 6987
rect 7849 6885 7883 6919
rect 9689 6817 9723 6851
rect 10333 6817 10367 6851
rect 46305 6817 46339 6851
rect 1961 6749 1995 6783
rect 3065 6749 3099 6783
rect 3893 6749 3927 6783
rect 4721 6749 4755 6783
rect 5181 6749 5215 6783
rect 8953 6749 8987 6783
rect 9597 6749 9631 6783
rect 9781 6749 9815 6783
rect 13093 6749 13127 6783
rect 7573 6681 7607 6715
rect 10609 6681 10643 6715
rect 46489 6681 46523 6715
rect 48145 6681 48179 6715
rect 2053 6613 2087 6647
rect 3157 6613 3191 6647
rect 3985 6613 4019 6647
rect 6929 6613 6963 6647
rect 8033 6613 8067 6647
rect 9045 6613 9079 6647
rect 12081 6613 12115 6647
rect 13185 6613 13219 6647
rect 12449 6409 12483 6443
rect 5365 6341 5399 6375
rect 9413 6341 9447 6375
rect 13277 6341 13311 6375
rect 1961 6273 1995 6307
rect 2605 6273 2639 6307
rect 4077 6273 4111 6307
rect 4721 6273 4755 6307
rect 5181 6273 5215 6307
rect 6377 6273 6411 6307
rect 8585 6273 8619 6307
rect 9597 6273 9631 6307
rect 9689 6273 9723 6307
rect 10333 6273 10367 6307
rect 12357 6273 12391 6307
rect 13093 6273 13127 6307
rect 13737 6273 13771 6307
rect 14381 6273 14415 6307
rect 45201 6273 45235 6307
rect 6653 6205 6687 6239
rect 10425 6205 10459 6239
rect 10701 6205 10735 6239
rect 45385 6205 45419 6239
rect 47041 6205 47075 6239
rect 4537 6137 4571 6171
rect 9413 6137 9447 6171
rect 14473 6137 14507 6171
rect 2053 6069 2087 6103
rect 2697 6069 2731 6103
rect 3433 6069 3467 6103
rect 3893 6069 3927 6103
rect 5549 6069 5583 6103
rect 8125 6069 8159 6103
rect 8677 6069 8711 6103
rect 13829 6069 13863 6103
rect 47777 6069 47811 6103
rect 3893 5865 3927 5899
rect 11621 5865 11655 5899
rect 11805 5865 11839 5899
rect 12449 5865 12483 5899
rect 9505 5797 9539 5831
rect 1961 5729 1995 5763
rect 9045 5729 9079 5763
rect 10701 5729 10735 5763
rect 10977 5729 11011 5763
rect 15025 5729 15059 5763
rect 31033 5729 31067 5763
rect 44465 5729 44499 5763
rect 46305 5729 46339 5763
rect 47133 5729 47167 5763
rect 2421 5661 2455 5695
rect 3065 5661 3099 5695
rect 3801 5661 3835 5695
rect 4445 5661 4479 5695
rect 6653 5661 6687 5695
rect 9137 5661 9171 5695
rect 10609 5661 10643 5695
rect 12265 5661 12299 5695
rect 13369 5661 13403 5695
rect 14289 5661 14323 5695
rect 14933 5661 14967 5695
rect 31677 5661 31711 5695
rect 32321 5661 32355 5695
rect 36369 5661 36403 5695
rect 37013 5661 37047 5695
rect 38393 5661 38427 5695
rect 40233 5661 40267 5695
rect 41613 5661 41647 5695
rect 43361 5661 43395 5695
rect 45017 5661 45051 5695
rect 45661 5661 45695 5695
rect 3157 5593 3191 5627
rect 4721 5593 4755 5627
rect 6929 5593 6963 5627
rect 11437 5593 11471 5627
rect 13461 5593 13495 5627
rect 45753 5593 45787 5627
rect 46489 5593 46523 5627
rect 2513 5525 2547 5559
rect 6193 5525 6227 5559
rect 8401 5525 8435 5559
rect 11637 5525 11671 5559
rect 14381 5525 14415 5559
rect 43453 5525 43487 5559
rect 45109 5525 45143 5559
rect 3617 5321 3651 5355
rect 4813 5321 4847 5355
rect 7021 5321 7055 5355
rect 7205 5321 7239 5355
rect 7389 5321 7423 5355
rect 10425 5321 10459 5355
rect 10517 5321 10551 5355
rect 10701 5321 10735 5355
rect 13277 5321 13311 5355
rect 2421 5253 2455 5287
rect 7113 5253 7147 5287
rect 8125 5253 8159 5287
rect 11805 5253 11839 5287
rect 2237 5185 2271 5219
rect 2973 5185 3007 5219
rect 3801 5185 3835 5219
rect 4445 5185 4479 5219
rect 5457 5185 5491 5219
rect 5641 5185 5675 5219
rect 6837 5185 6871 5219
rect 10333 5185 10367 5219
rect 16681 5185 16715 5219
rect 17325 5185 17359 5219
rect 18337 5185 18371 5219
rect 20269 5185 20303 5219
rect 21833 5185 21867 5219
rect 28365 5185 28399 5219
rect 29009 5185 29043 5219
rect 30481 5185 30515 5219
rect 31125 5185 31159 5219
rect 32137 5185 32171 5219
rect 32781 5185 32815 5219
rect 33425 5185 33459 5219
rect 34069 5185 34103 5219
rect 35357 5185 35391 5219
rect 37289 5185 37323 5219
rect 37933 5185 37967 5219
rect 38577 5185 38611 5219
rect 40509 5185 40543 5219
rect 41153 5185 41187 5219
rect 42441 5185 42475 5219
rect 43729 5185 43763 5219
rect 44373 5185 44407 5219
rect 45201 5185 45235 5219
rect 47593 5185 47627 5219
rect 4353 5117 4387 5151
rect 5549 5117 5583 5151
rect 5733 5117 5767 5151
rect 7849 5117 7883 5151
rect 11529 5117 11563 5151
rect 45385 5117 45419 5151
rect 47041 5117 47075 5151
rect 1685 5049 1719 5083
rect 5273 5049 5307 5083
rect 10149 5049 10183 5083
rect 15117 5049 15151 5083
rect 30573 5049 30607 5083
rect 33517 5049 33551 5083
rect 36185 5049 36219 5083
rect 3065 4981 3099 5015
rect 9597 4981 9631 5015
rect 14381 4981 14415 5015
rect 15761 4981 15795 5015
rect 16773 4981 16807 5015
rect 17417 4981 17451 5015
rect 18429 4981 18463 5015
rect 19165 4981 19199 5015
rect 19809 4981 19843 5015
rect 20361 4981 20395 5015
rect 21281 4981 21315 5015
rect 21925 4981 21959 5015
rect 23213 4981 23247 5015
rect 24133 4981 24167 5015
rect 24777 4981 24811 5015
rect 28457 4981 28491 5015
rect 29101 4981 29135 5015
rect 31217 4981 31251 5015
rect 32229 4981 32263 5015
rect 32873 4981 32907 5015
rect 34161 4981 34195 5015
rect 34897 4981 34931 5015
rect 35449 4981 35483 5015
rect 37381 4981 37415 5015
rect 38025 4981 38059 5015
rect 38669 4981 38703 5015
rect 39405 4981 39439 5015
rect 40049 4981 40083 5015
rect 40601 4981 40635 5015
rect 41245 4981 41279 5015
rect 42533 4981 42567 5015
rect 43269 4981 43303 5015
rect 43821 4981 43855 5015
rect 44465 4981 44499 5015
rect 47685 4981 47719 5015
rect 3249 4777 3283 4811
rect 32137 4777 32171 4811
rect 33241 4777 33275 4811
rect 44373 4777 44407 4811
rect 14749 4709 14783 4743
rect 19809 4709 19843 4743
rect 1685 4641 1719 4675
rect 2881 4641 2915 4675
rect 3801 4641 3835 4675
rect 4261 4641 4295 4675
rect 6285 4641 6319 4675
rect 6469 4641 6503 4675
rect 6929 4641 6963 4675
rect 8953 4641 8987 4675
rect 9137 4641 9171 4675
rect 9781 4641 9815 4675
rect 11437 4641 11471 4675
rect 27353 4641 27387 4675
rect 45845 4641 45879 4675
rect 46029 4641 46063 4675
rect 46489 4641 46523 4675
rect 1593 4573 1627 4607
rect 1777 4573 1811 4607
rect 2237 4573 2271 4607
rect 3065 4573 3099 4607
rect 15301 4573 15335 4607
rect 16129 4573 16163 4607
rect 16773 4573 16807 4607
rect 17417 4573 17451 4607
rect 18061 4573 18095 4607
rect 18521 4573 18555 4607
rect 20269 4573 20303 4607
rect 20545 4573 20579 4607
rect 21925 4573 21959 4607
rect 22385 4573 22419 4607
rect 23029 4573 23063 4607
rect 23673 4573 23707 4607
rect 24593 4573 24627 4607
rect 25237 4573 25271 4607
rect 26065 4573 26099 4607
rect 28089 4573 28123 4607
rect 28549 4573 28583 4607
rect 29745 4573 29779 4607
rect 30389 4573 30423 4607
rect 31033 4573 31067 4607
rect 33977 4573 34011 4607
rect 34897 4573 34931 4607
rect 35357 4573 35391 4607
rect 36185 4573 36219 4607
rect 36645 4573 36679 4607
rect 37749 4573 37783 4607
rect 38209 4573 38243 4607
rect 39037 4573 39071 4607
rect 39865 4573 39899 4607
rect 40785 4573 40819 4607
rect 40969 4573 41003 4607
rect 41429 4573 41463 4607
rect 42257 4573 42291 4607
rect 42717 4573 42751 4607
rect 43545 4573 43579 4607
rect 44281 4573 44315 4607
rect 45201 4573 45235 4607
rect 3985 4505 4019 4539
rect 11621 4505 11655 4539
rect 13277 4505 13311 4539
rect 14565 4505 14599 4539
rect 19625 4505 19659 4539
rect 27905 4505 27939 4539
rect 32045 4505 32079 4539
rect 33149 4505 33183 4539
rect 37565 4505 37599 4539
rect 45385 4505 45419 4539
rect 2329 4437 2363 4471
rect 15393 4437 15427 4471
rect 18613 4437 18647 4471
rect 22477 4437 22511 4471
rect 23121 4437 23155 4471
rect 23765 4437 23799 4471
rect 24685 4437 24719 4471
rect 25329 4437 25363 4471
rect 28641 4437 28675 4471
rect 35449 4437 35483 4471
rect 36737 4437 36771 4471
rect 38301 4437 38335 4471
rect 39957 4437 39991 4471
rect 41521 4437 41555 4471
rect 42809 4437 42843 4471
rect 23305 4233 23339 4267
rect 15669 4165 15703 4199
rect 18705 4165 18739 4199
rect 20913 4165 20947 4199
rect 21097 4165 21131 4199
rect 24041 4165 24075 4199
rect 28457 4165 28491 4199
rect 32321 4165 32355 4199
rect 34897 4165 34931 4199
rect 37565 4165 37599 4199
rect 1593 4097 1627 4131
rect 3985 4097 4019 4131
rect 12541 4097 12575 4131
rect 15853 4097 15887 4131
rect 17233 4097 17267 4131
rect 17877 4097 17911 4131
rect 18521 4097 18555 4131
rect 22477 4097 22511 4131
rect 23213 4097 23247 4131
rect 23857 4097 23891 4131
rect 27629 4097 27663 4131
rect 31217 4097 31251 4131
rect 32137 4097 32171 4131
rect 42625 4097 42659 4131
rect 1777 4029 1811 4063
rect 2053 4029 2087 4063
rect 4169 4029 4203 4063
rect 4445 4029 4479 4063
rect 6837 4029 6871 4063
rect 7021 4029 7055 4063
rect 7297 4029 7331 4063
rect 9137 4029 9171 4063
rect 9321 4029 9355 4063
rect 10977 4029 11011 4063
rect 12817 4029 12851 4063
rect 13093 4029 13127 4063
rect 13277 4029 13311 4063
rect 13461 4029 13495 4063
rect 15117 4029 15151 4063
rect 20085 4029 20119 4063
rect 24501 4029 24535 4063
rect 28273 4029 28307 4063
rect 29837 4029 29871 4063
rect 32965 4029 32999 4063
rect 34713 4029 34747 4063
rect 36277 4029 36311 4063
rect 37381 4029 37415 4063
rect 38117 4029 38151 4063
rect 40049 4029 40083 4063
rect 40233 4029 40267 4063
rect 41613 4029 41647 4063
rect 42809 4029 42843 4063
rect 44005 4029 44039 4063
rect 45017 4029 45051 4063
rect 45201 4029 45235 4063
rect 45845 4029 45879 4063
rect 47777 3961 47811 3995
rect 17325 3893 17359 3927
rect 17969 3893 18003 3927
rect 22017 3893 22051 3927
rect 22569 3893 22603 3927
rect 26341 3893 26375 3927
rect 27169 3893 27203 3927
rect 27721 3893 27755 3927
rect 30757 3893 30791 3927
rect 31309 3893 31343 3927
rect 47501 3621 47535 3655
rect 1409 3553 1443 3587
rect 1869 3553 1903 3587
rect 4261 3553 4295 3587
rect 4445 3553 4479 3587
rect 5917 3553 5951 3587
rect 6561 3553 6595 3587
rect 8953 3553 8987 3587
rect 10425 3553 10459 3587
rect 11253 3553 11287 3587
rect 14197 3553 14231 3587
rect 16497 3553 16531 3587
rect 16681 3553 16715 3587
rect 18153 3553 18187 3587
rect 19257 3553 19291 3587
rect 19441 3553 19475 3587
rect 20729 3553 20763 3587
rect 21649 3553 21683 3587
rect 26525 3553 26559 3587
rect 29561 3553 29595 3587
rect 29745 3553 29779 3587
rect 31861 3553 31895 3587
rect 32045 3553 32079 3587
rect 32321 3553 32355 3587
rect 34713 3553 34747 3587
rect 35173 3553 35207 3587
rect 37013 3553 37047 3587
rect 37197 3553 37231 3587
rect 37473 3553 37507 3587
rect 39865 3553 39899 3587
rect 40325 3553 40359 3587
rect 42165 3553 42199 3587
rect 42349 3553 42383 3587
rect 42901 3553 42935 3587
rect 45201 3553 45235 3587
rect 48053 3553 48087 3587
rect 24961 3485 24995 3519
rect 25697 3485 25731 3519
rect 27997 3485 28031 3519
rect 28825 3485 28859 3519
rect 45017 3485 45051 3519
rect 47961 3485 47995 3519
rect 1593 3417 1627 3451
rect 6745 3417 6779 3451
rect 8401 3417 8435 3451
rect 9137 3417 9171 3451
rect 11437 3417 11471 3451
rect 13093 3417 13127 3451
rect 14381 3417 14415 3451
rect 16037 3417 16071 3451
rect 21833 3417 21867 3451
rect 23489 3417 23523 3451
rect 25881 3417 25915 3451
rect 31401 3417 31435 3451
rect 34897 3417 34931 3451
rect 40049 3417 40083 3451
rect 46857 3417 46891 3451
rect 25053 3349 25087 3383
rect 28089 3349 28123 3383
rect 1869 3077 1903 3111
rect 4169 3077 4203 3111
rect 7021 3077 7055 3111
rect 10977 3077 11011 3111
rect 14473 3077 14507 3111
rect 18981 3077 19015 3111
rect 19625 3077 19659 3111
rect 22477 3077 22511 3111
rect 24777 3077 24811 3111
rect 27169 3077 27203 3111
rect 29469 3077 29503 3111
rect 32321 3077 32355 3111
rect 34621 3077 34655 3111
rect 37473 3077 37507 3111
rect 39773 3077 39807 3111
rect 42625 3077 42659 3111
rect 44925 3077 44959 3111
rect 1685 3009 1719 3043
rect 6837 3009 6871 3043
rect 16129 3009 16163 3043
rect 17141 3009 17175 3043
rect 22293 3009 22327 3043
rect 26985 3009 27019 3043
rect 29285 3009 29319 3043
rect 32137 3009 32171 3043
rect 34437 3009 34471 3043
rect 39589 3009 39623 3043
rect 42441 3009 42475 3043
rect 47777 3009 47811 3043
rect 2697 2941 2731 2975
rect 3985 2941 4019 2975
rect 5365 2941 5399 2975
rect 8677 2941 8711 2975
rect 9137 2941 9171 2975
rect 9321 2941 9355 2975
rect 11989 2941 12023 2975
rect 12173 2941 12207 2975
rect 13829 2941 13863 2975
rect 14289 2941 14323 2975
rect 17325 2941 17359 2975
rect 19441 2941 19475 2975
rect 21281 2941 21315 2975
rect 23949 2941 23983 2975
rect 24593 2941 24627 2975
rect 25973 2941 26007 2975
rect 27445 2941 27479 2975
rect 29745 2941 29779 2975
rect 32597 2941 32631 2975
rect 34897 2941 34931 2975
rect 37289 2941 37323 2975
rect 37749 2941 37783 2975
rect 40049 2941 40083 2975
rect 42901 2941 42935 2975
rect 44741 2941 44775 2975
rect 45201 2941 45235 2975
rect 47777 2601 47811 2635
rect 1409 2465 1443 2499
rect 1593 2465 1627 2499
rect 2053 2465 2087 2499
rect 3985 2465 4019 2499
rect 4169 2465 4203 2499
rect 4629 2465 4663 2499
rect 6561 2465 6595 2499
rect 7757 2465 7791 2499
rect 8953 2465 8987 2499
rect 9413 2465 9447 2499
rect 11621 2465 11655 2499
rect 16865 2465 16899 2499
rect 17049 2465 17083 2499
rect 19441 2465 19475 2499
rect 19625 2465 19659 2499
rect 22017 2465 22051 2499
rect 22201 2465 22235 2499
rect 23489 2465 23523 2499
rect 24593 2465 24627 2499
rect 24777 2465 24811 2499
rect 25237 2465 25271 2499
rect 26985 2465 27019 2499
rect 27169 2465 27203 2499
rect 27813 2465 27847 2499
rect 29561 2465 29595 2499
rect 30941 2465 30975 2499
rect 32137 2465 32171 2499
rect 32321 2465 32355 2499
rect 32597 2465 32631 2499
rect 35173 2465 35207 2499
rect 37289 2465 37323 2499
rect 37473 2465 37507 2499
rect 38393 2465 38427 2499
rect 39865 2465 39899 2499
rect 40049 2465 40083 2499
rect 40325 2465 40359 2499
rect 42441 2465 42475 2499
rect 42625 2465 42659 2499
rect 42901 2465 42935 2499
rect 45017 2465 45051 2499
rect 45661 2465 45695 2499
rect 14289 2397 14323 2431
rect 34713 2397 34747 2431
rect 6745 2329 6779 2363
rect 9137 2329 9171 2363
rect 11805 2329 11839 2363
rect 13461 2329 13495 2363
rect 14473 2329 14507 2363
rect 16129 2329 16163 2363
rect 18705 2329 18739 2363
rect 21281 2329 21315 2363
rect 29745 2329 29779 2363
rect 34897 2329 34931 2363
rect 45201 2329 45235 2363
<< metal1 >>
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 2041 47175 2099 47181
rect 2041 47141 2053 47175
rect 2087 47172 2099 47175
rect 2222 47172 2228 47184
rect 2087 47144 2228 47172
rect 2087 47141 2099 47144
rect 2041 47135 2099 47141
rect 2222 47132 2228 47144
rect 2280 47132 2286 47184
rect 34882 47132 34888 47184
rect 34940 47172 34946 47184
rect 35161 47175 35219 47181
rect 35161 47172 35173 47175
rect 34940 47144 35173 47172
rect 34940 47132 34946 47144
rect 35161 47141 35173 47144
rect 35207 47141 35219 47175
rect 35161 47135 35219 47141
rect 1762 46996 1768 47048
rect 1820 47036 1826 47048
rect 1857 47039 1915 47045
rect 1857 47036 1869 47039
rect 1820 47008 1869 47036
rect 1820 46996 1826 47008
rect 1857 47005 1869 47008
rect 1903 47005 1915 47039
rect 5258 47036 5264 47048
rect 5219 47008 5264 47036
rect 1857 46999 1915 47005
rect 5258 46996 5264 47008
rect 5316 46996 5322 47048
rect 21818 47036 21824 47048
rect 21779 47008 21824 47036
rect 21818 46996 21824 47008
rect 21876 46996 21882 47048
rect 24946 46996 24952 47048
rect 25004 47036 25010 47048
rect 25041 47039 25099 47045
rect 25041 47036 25053 47039
rect 25004 47008 25053 47036
rect 25004 46996 25010 47008
rect 25041 47005 25053 47008
rect 25087 47005 25099 47039
rect 25041 46999 25099 47005
rect 28258 46996 28264 47048
rect 28316 47036 28322 47048
rect 28353 47039 28411 47045
rect 28353 47036 28365 47039
rect 28316 47008 28365 47036
rect 28316 46996 28322 47008
rect 28353 47005 28365 47008
rect 28399 47005 28411 47039
rect 28353 46999 28411 47005
rect 31754 46996 31760 47048
rect 31812 47036 31818 47048
rect 32125 47039 32183 47045
rect 32125 47036 32137 47039
rect 31812 47008 32137 47036
rect 31812 46996 31818 47008
rect 32125 47005 32137 47008
rect 32171 47005 32183 47039
rect 32125 46999 32183 47005
rect 34790 46996 34796 47048
rect 34848 47036 34854 47048
rect 34977 47039 35035 47045
rect 34977 47036 34989 47039
rect 34848 47008 34989 47036
rect 34848 46996 34854 47008
rect 34977 47005 34989 47008
rect 35023 47005 35035 47039
rect 34977 46999 35035 47005
rect 38194 46996 38200 47048
rect 38252 47036 38258 47048
rect 38289 47039 38347 47045
rect 38289 47036 38301 47039
rect 38252 47008 38301 47036
rect 38252 46996 38258 47008
rect 38289 47005 38301 47008
rect 38335 47005 38347 47039
rect 38289 46999 38347 47005
rect 44818 46996 44824 47048
rect 44876 47036 44882 47048
rect 45465 47039 45523 47045
rect 45465 47036 45477 47039
rect 44876 47008 45477 47036
rect 44876 46996 44882 47008
rect 45465 47005 45477 47008
rect 45511 47005 45523 47039
rect 45465 46999 45523 47005
rect 47673 47039 47731 47045
rect 47673 47005 47685 47039
rect 47719 47036 47731 47039
rect 48130 47036 48136 47048
rect 47719 47008 48136 47036
rect 47719 47005 47731 47008
rect 47673 46999 47731 47005
rect 48130 46996 48136 47008
rect 48188 46996 48194 47048
rect 5629 46971 5687 46977
rect 5629 46937 5641 46971
rect 5675 46968 5687 46971
rect 8202 46968 8208 46980
rect 5675 46940 8208 46968
rect 5675 46937 5687 46940
rect 5629 46931 5687 46937
rect 8202 46928 8208 46940
rect 8260 46928 8266 46980
rect 42889 46971 42947 46977
rect 42889 46968 42901 46971
rect 42812 46940 42901 46968
rect 22002 46900 22008 46912
rect 21963 46872 22008 46900
rect 22002 46860 22008 46872
rect 22060 46860 22066 46912
rect 25222 46900 25228 46912
rect 25183 46872 25228 46900
rect 25222 46860 25228 46872
rect 25280 46860 25286 46912
rect 28534 46900 28540 46912
rect 28495 46872 28540 46900
rect 28534 46860 28540 46872
rect 28592 46860 28598 46912
rect 32306 46900 32312 46912
rect 32267 46872 32312 46900
rect 32306 46860 32312 46872
rect 32364 46860 32370 46912
rect 38470 46900 38476 46912
rect 38431 46872 38476 46900
rect 38470 46860 38476 46872
rect 38528 46860 38534 46912
rect 41506 46860 41512 46912
rect 41564 46900 41570 46912
rect 42812 46900 42840 46940
rect 42889 46937 42901 46940
rect 42935 46937 42947 46971
rect 47946 46968 47952 46980
rect 47907 46940 47952 46968
rect 42889 46931 42947 46937
rect 47946 46928 47952 46940
rect 48004 46928 48010 46980
rect 42978 46900 42984 46912
rect 41564 46872 42840 46900
rect 42939 46872 42984 46900
rect 41564 46860 41570 46872
rect 42978 46860 42984 46872
rect 43036 46860 43042 46912
rect 45554 46860 45560 46912
rect 45612 46900 45618 46912
rect 45612 46872 45657 46900
rect 45612 46860 45618 46872
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 10318 8956 10324 8968
rect 10279 8928 10324 8956
rect 10318 8916 10324 8928
rect 10376 8956 10382 8968
rect 12526 8956 12532 8968
rect 10376 8928 12532 8956
rect 10376 8916 10382 8928
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 10410 8820 10416 8832
rect 10371 8792 10416 8820
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 11882 8780 11888 8832
rect 11940 8820 11946 8832
rect 12621 8823 12679 8829
rect 12621 8820 12633 8823
rect 11940 8792 12633 8820
rect 11940 8780 11946 8792
rect 12621 8789 12633 8792
rect 12667 8789 12679 8823
rect 12621 8783 12679 8789
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 7650 8480 7656 8492
rect 7611 8452 7656 8480
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8449 8447 8483
rect 8389 8443 8447 8449
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8480 9091 8483
rect 9677 8483 9735 8489
rect 9677 8480 9689 8483
rect 9079 8452 9689 8480
rect 9079 8449 9091 8452
rect 9033 8443 9091 8449
rect 9677 8449 9689 8452
rect 9723 8480 9735 8483
rect 10962 8480 10968 8492
rect 9723 8452 10968 8480
rect 9723 8449 9735 8452
rect 9677 8443 9735 8449
rect 8404 8412 8432 8443
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 47578 8440 47584 8492
rect 47636 8480 47642 8492
rect 47857 8483 47915 8489
rect 47857 8480 47869 8483
rect 47636 8452 47869 8480
rect 47636 8440 47642 8452
rect 47857 8449 47869 8452
rect 47903 8449 47915 8483
rect 47857 8443 47915 8449
rect 9582 8412 9588 8424
rect 8404 8384 9588 8412
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 1578 8304 1584 8356
rect 1636 8344 1642 8356
rect 1857 8347 1915 8353
rect 1857 8344 1869 8347
rect 1636 8316 1869 8344
rect 1636 8304 1642 8316
rect 1857 8313 1869 8316
rect 1903 8313 1915 8347
rect 7742 8344 7748 8356
rect 7703 8316 7748 8344
rect 1857 8307 1915 8313
rect 7742 8304 7748 8316
rect 7800 8304 7806 8356
rect 8481 8347 8539 8353
rect 8481 8313 8493 8347
rect 8527 8344 8539 8347
rect 8846 8344 8852 8356
rect 8527 8316 8852 8344
rect 8527 8313 8539 8316
rect 8481 8307 8539 8313
rect 8846 8304 8852 8316
rect 8904 8304 8910 8356
rect 9030 8304 9036 8356
rect 9088 8344 9094 8356
rect 9125 8347 9183 8353
rect 9125 8344 9137 8347
rect 9088 8316 9137 8344
rect 9088 8304 9094 8316
rect 9125 8313 9137 8316
rect 9171 8313 9183 8347
rect 9125 8307 9183 8313
rect 9306 8304 9312 8356
rect 9364 8344 9370 8356
rect 9769 8347 9827 8353
rect 9769 8344 9781 8347
rect 9364 8316 9781 8344
rect 9364 8304 9370 8316
rect 9769 8313 9781 8316
rect 9815 8313 9827 8347
rect 9769 8307 9827 8313
rect 45370 8304 45376 8356
rect 45428 8344 45434 8356
rect 47949 8347 48007 8353
rect 47949 8344 47961 8347
rect 45428 8316 47961 8344
rect 45428 8304 45434 8316
rect 47949 8313 47961 8316
rect 47995 8313 48007 8347
rect 47949 8307 48007 8313
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 8478 8032 8484 8084
rect 8536 8072 8542 8084
rect 10321 8075 10379 8081
rect 10321 8072 10333 8075
rect 8536 8044 10333 8072
rect 8536 8032 8542 8044
rect 10321 8041 10333 8044
rect 10367 8041 10379 8075
rect 10321 8035 10379 8041
rect 1394 7896 1400 7948
rect 1452 7936 1458 7948
rect 2593 7939 2651 7945
rect 2593 7936 2605 7939
rect 1452 7908 2605 7936
rect 1452 7896 1458 7908
rect 2593 7905 2605 7908
rect 2639 7905 2651 7939
rect 10318 7936 10324 7948
rect 2593 7899 2651 7905
rect 8220 7908 10324 7936
rect 8220 7880 8248 7908
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 1854 7868 1860 7880
rect 1815 7840 1860 7868
rect 1854 7828 1860 7840
rect 1912 7828 1918 7880
rect 6086 7868 6092 7880
rect 6047 7840 6092 7868
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7837 7067 7871
rect 8202 7868 8208 7880
rect 8163 7840 8208 7868
rect 7009 7831 7067 7837
rect 7024 7800 7052 7831
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 9582 7868 9588 7880
rect 9447 7840 9588 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 10505 7871 10563 7877
rect 10505 7837 10517 7871
rect 10551 7837 10563 7871
rect 10962 7868 10968 7880
rect 10923 7840 10968 7868
rect 10505 7831 10563 7837
rect 7190 7800 7196 7812
rect 7024 7772 7196 7800
rect 7190 7760 7196 7772
rect 7248 7800 7254 7812
rect 7650 7800 7656 7812
rect 7248 7772 7656 7800
rect 7248 7760 7254 7772
rect 7650 7760 7656 7772
rect 7708 7800 7714 7812
rect 8389 7803 8447 7809
rect 8389 7800 8401 7803
rect 7708 7772 8401 7800
rect 7708 7760 7714 7772
rect 8389 7769 8401 7772
rect 8435 7800 8447 7803
rect 8938 7800 8944 7812
rect 8435 7772 8944 7800
rect 8435 7769 8447 7772
rect 8389 7763 8447 7769
rect 8938 7760 8944 7772
rect 8996 7760 9002 7812
rect 10045 7803 10103 7809
rect 10045 7769 10057 7803
rect 10091 7800 10103 7803
rect 10226 7800 10232 7812
rect 10091 7772 10232 7800
rect 10091 7769 10103 7772
rect 10045 7763 10103 7769
rect 10226 7760 10232 7772
rect 10284 7800 10290 7812
rect 10520 7800 10548 7831
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 47118 7868 47124 7880
rect 47079 7840 47124 7868
rect 47118 7828 47124 7840
rect 47176 7828 47182 7880
rect 47578 7868 47584 7880
rect 47539 7840 47584 7868
rect 47578 7828 47584 7840
rect 47636 7828 47642 7880
rect 47946 7800 47952 7812
rect 10284 7772 47952 7800
rect 10284 7760 10290 7772
rect 47946 7760 47952 7772
rect 48004 7760 48010 7812
rect 5166 7692 5172 7744
rect 5224 7732 5230 7744
rect 6181 7735 6239 7741
rect 6181 7732 6193 7735
rect 5224 7704 6193 7732
rect 5224 7692 5230 7704
rect 6181 7701 6193 7704
rect 6227 7701 6239 7735
rect 7098 7732 7104 7744
rect 7059 7704 7104 7732
rect 6181 7695 6239 7701
rect 7098 7692 7104 7704
rect 7156 7692 7162 7744
rect 9214 7692 9220 7744
rect 9272 7732 9278 7744
rect 9493 7735 9551 7741
rect 9493 7732 9505 7735
rect 9272 7704 9505 7732
rect 9272 7692 9278 7704
rect 9493 7701 9505 7704
rect 9539 7701 9551 7735
rect 11054 7732 11060 7744
rect 11015 7704 11060 7732
rect 9493 7695 9551 7701
rect 11054 7692 11060 7704
rect 11112 7692 11118 7744
rect 47670 7732 47676 7744
rect 47631 7704 47676 7732
rect 47670 7692 47676 7704
rect 47728 7692 47734 7744
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 8478 7460 8484 7472
rect 6748 7432 8484 7460
rect 1946 7392 1952 7404
rect 1907 7364 1952 7392
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 4982 7392 4988 7404
rect 4943 7364 4988 7392
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 5592 7364 5641 7392
rect 5592 7352 5598 7364
rect 5629 7361 5641 7364
rect 5675 7392 5687 7395
rect 6086 7392 6092 7404
rect 5675 7364 6092 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 6086 7352 6092 7364
rect 6144 7392 6150 7404
rect 6638 7392 6644 7404
rect 6144 7364 6644 7392
rect 6144 7352 6150 7364
rect 6638 7352 6644 7364
rect 6696 7352 6702 7404
rect 6748 7401 6776 7432
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7361 6791 7395
rect 7190 7392 7196 7404
rect 7151 7364 7196 7392
rect 6733 7355 6791 7361
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 7944 7401 7972 7432
rect 8478 7420 8484 7432
rect 8536 7420 8542 7472
rect 10410 7460 10416 7472
rect 9430 7432 10416 7460
rect 10410 7420 10416 7432
rect 10468 7420 10474 7472
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 10689 7395 10747 7401
rect 10689 7361 10701 7395
rect 10735 7392 10747 7395
rect 10962 7392 10968 7404
rect 10735 7364 10968 7392
rect 10735 7361 10747 7364
rect 10689 7355 10747 7361
rect 10962 7352 10968 7364
rect 11020 7392 11026 7404
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 11020 7364 11529 7392
rect 11020 7352 11026 7364
rect 11517 7361 11529 7364
rect 11563 7392 11575 7395
rect 12434 7392 12440 7404
rect 11563 7364 12440 7392
rect 11563 7361 11575 7364
rect 11517 7355 11575 7361
rect 12434 7352 12440 7364
rect 12492 7352 12498 7404
rect 47578 7392 47584 7404
rect 47539 7364 47584 7392
rect 47578 7352 47584 7364
rect 47636 7352 47642 7404
rect 8205 7327 8263 7333
rect 8205 7293 8217 7327
rect 8251 7324 8263 7327
rect 9490 7324 9496 7336
rect 8251 7296 9496 7324
rect 8251 7293 8263 7296
rect 8205 7287 8263 7293
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 45278 7284 45284 7336
rect 45336 7324 45342 7336
rect 47673 7327 47731 7333
rect 47673 7324 47685 7327
rect 45336 7296 47685 7324
rect 45336 7284 45342 7296
rect 47673 7293 47685 7296
rect 47719 7293 47731 7327
rect 47673 7287 47731 7293
rect 6362 7216 6368 7268
rect 6420 7256 6426 7268
rect 6549 7259 6607 7265
rect 6549 7256 6561 7259
rect 6420 7228 6561 7256
rect 6420 7216 6426 7228
rect 6549 7225 6561 7228
rect 6595 7225 6607 7259
rect 6549 7219 6607 7225
rect 11146 7216 11152 7268
rect 11204 7256 11210 7268
rect 11609 7259 11667 7265
rect 11609 7256 11621 7259
rect 11204 7228 11621 7256
rect 11204 7216 11210 7228
rect 11609 7225 11621 7228
rect 11655 7225 11667 7259
rect 11609 7219 11667 7225
rect 45462 7216 45468 7268
rect 45520 7256 45526 7268
rect 47029 7259 47087 7265
rect 47029 7256 47041 7259
rect 45520 7228 47041 7256
rect 45520 7216 45526 7228
rect 47029 7225 47041 7228
rect 47075 7225 47087 7259
rect 47029 7219 47087 7225
rect 1762 7148 1768 7200
rect 1820 7188 1826 7200
rect 2041 7191 2099 7197
rect 2041 7188 2053 7191
rect 1820 7160 2053 7188
rect 1820 7148 1826 7160
rect 2041 7157 2053 7160
rect 2087 7157 2099 7191
rect 2041 7151 2099 7157
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 3329 7191 3387 7197
rect 3329 7188 3341 7191
rect 2832 7160 3341 7188
rect 2832 7148 2838 7160
rect 3329 7157 3341 7160
rect 3375 7157 3387 7191
rect 5074 7188 5080 7200
rect 5035 7160 5080 7188
rect 3329 7151 3387 7157
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 5721 7191 5779 7197
rect 5721 7157 5733 7191
rect 5767 7188 5779 7191
rect 6454 7188 6460 7200
rect 5767 7160 6460 7188
rect 5767 7157 5779 7160
rect 5721 7151 5779 7157
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 7282 7188 7288 7200
rect 7243 7160 7288 7188
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 9677 7191 9735 7197
rect 9677 7157 9689 7191
rect 9723 7188 9735 7191
rect 9858 7188 9864 7200
rect 9723 7160 9864 7188
rect 9723 7157 9735 7160
rect 9677 7151 9735 7157
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 10781 7191 10839 7197
rect 10781 7157 10793 7191
rect 10827 7188 10839 7191
rect 11422 7188 11428 7200
rect 10827 7160 11428 7188
rect 10827 7157 10839 7160
rect 10781 7151 10839 7157
rect 11422 7148 11428 7160
rect 11480 7148 11486 7200
rect 46382 7188 46388 7200
rect 46343 7160 46388 7188
rect 46382 7148 46388 7160
rect 46440 7148 46446 7200
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 5074 6944 5080 6996
rect 5132 6984 5138 6996
rect 5426 6987 5484 6993
rect 5426 6984 5438 6987
rect 5132 6956 5438 6984
rect 5132 6944 5138 6956
rect 5426 6953 5438 6956
rect 5472 6953 5484 6987
rect 5426 6947 5484 6953
rect 7837 6919 7895 6925
rect 7837 6885 7849 6919
rect 7883 6885 7895 6919
rect 7837 6879 7895 6885
rect 5534 6848 5540 6860
rect 3896 6820 5540 6848
rect 1946 6780 1952 6792
rect 1907 6752 1952 6780
rect 1946 6740 1952 6752
rect 2004 6780 2010 6792
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 2004 6752 3065 6780
rect 2004 6740 2010 6752
rect 3053 6749 3065 6752
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 3326 6740 3332 6792
rect 3384 6780 3390 6792
rect 3896 6789 3924 6820
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 5810 6808 5816 6860
rect 5868 6848 5874 6860
rect 7852 6848 7880 6879
rect 5868 6820 7880 6848
rect 5868 6808 5874 6820
rect 9490 6808 9496 6860
rect 9548 6848 9554 6860
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 9548 6820 9689 6848
rect 9548 6808 9554 6820
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 10226 6808 10232 6860
rect 10284 6848 10290 6860
rect 10321 6851 10379 6857
rect 10321 6848 10333 6851
rect 10284 6820 10333 6848
rect 10284 6808 10290 6820
rect 10321 6817 10333 6820
rect 10367 6817 10379 6851
rect 10321 6811 10379 6817
rect 46293 6851 46351 6857
rect 46293 6817 46305 6851
rect 46339 6848 46351 6851
rect 47118 6848 47124 6860
rect 46339 6820 47124 6848
rect 46339 6817 46351 6820
rect 46293 6811 46351 6817
rect 47118 6808 47124 6820
rect 47176 6808 47182 6860
rect 3881 6783 3939 6789
rect 3881 6780 3893 6783
rect 3384 6752 3893 6780
rect 3384 6740 3390 6752
rect 3881 6749 3893 6752
rect 3927 6749 3939 6783
rect 3881 6743 3939 6749
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 4798 6780 4804 6792
rect 4755 6752 4804 6780
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 4798 6740 4804 6752
rect 4856 6740 4862 6792
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6749 5227 6783
rect 8938 6780 8944 6792
rect 8899 6752 8944 6780
rect 5169 6743 5227 6749
rect 4614 6672 4620 6724
rect 4672 6712 4678 6724
rect 5184 6712 5212 6743
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 9585 6783 9643 6789
rect 9585 6780 9597 6783
rect 9456 6752 9597 6780
rect 9456 6740 9462 6752
rect 9585 6749 9597 6752
rect 9631 6749 9643 6783
rect 9766 6780 9772 6792
rect 9727 6752 9772 6780
rect 9585 6743 9643 6749
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 12526 6740 12532 6792
rect 12584 6780 12590 6792
rect 13081 6783 13139 6789
rect 13081 6780 13093 6783
rect 12584 6752 13093 6780
rect 12584 6740 12590 6752
rect 13081 6749 13093 6752
rect 13127 6749 13139 6783
rect 13081 6743 13139 6749
rect 5718 6712 5724 6724
rect 4672 6684 5724 6712
rect 4672 6672 4678 6684
rect 5718 6672 5724 6684
rect 5776 6672 5782 6724
rect 7098 6712 7104 6724
rect 6670 6684 7104 6712
rect 7098 6672 7104 6684
rect 7156 6672 7162 6724
rect 7558 6712 7564 6724
rect 7519 6684 7564 6712
rect 7558 6672 7564 6684
rect 7616 6672 7622 6724
rect 10594 6712 10600 6724
rect 10555 6684 10600 6712
rect 10594 6672 10600 6684
rect 10652 6672 10658 6724
rect 11882 6712 11888 6724
rect 11822 6684 11888 6712
rect 11882 6672 11888 6684
rect 11940 6672 11946 6724
rect 46477 6715 46535 6721
rect 46477 6681 46489 6715
rect 46523 6712 46535 6715
rect 47670 6712 47676 6724
rect 46523 6684 47676 6712
rect 46523 6681 46535 6684
rect 46477 6675 46535 6681
rect 47670 6672 47676 6684
rect 47728 6672 47734 6724
rect 48133 6715 48191 6721
rect 48133 6681 48145 6715
rect 48179 6712 48191 6715
rect 49050 6712 49056 6724
rect 48179 6684 49056 6712
rect 48179 6681 48191 6684
rect 48133 6675 48191 6681
rect 49050 6672 49056 6684
rect 49108 6672 49114 6724
rect 2038 6644 2044 6656
rect 1999 6616 2044 6644
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 3142 6644 3148 6656
rect 3103 6616 3148 6644
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 3973 6647 4031 6653
rect 3973 6613 3985 6647
rect 4019 6644 4031 6647
rect 4706 6644 4712 6656
rect 4019 6616 4712 6644
rect 4019 6613 4031 6616
rect 3973 6607 4031 6613
rect 4706 6604 4712 6616
rect 4764 6604 4770 6656
rect 4982 6604 4988 6656
rect 5040 6644 5046 6656
rect 5626 6644 5632 6656
rect 5040 6616 5632 6644
rect 5040 6604 5046 6616
rect 5626 6604 5632 6616
rect 5684 6644 5690 6656
rect 6917 6647 6975 6653
rect 6917 6644 6929 6647
rect 5684 6616 6929 6644
rect 5684 6604 5690 6616
rect 6917 6613 6929 6616
rect 6963 6613 6975 6647
rect 8018 6644 8024 6656
rect 7979 6616 8024 6644
rect 6917 6607 6975 6613
rect 8018 6604 8024 6616
rect 8076 6604 8082 6656
rect 9033 6647 9091 6653
rect 9033 6613 9045 6647
rect 9079 6644 9091 6647
rect 9122 6644 9128 6656
rect 9079 6616 9128 6644
rect 9079 6613 9091 6616
rect 9033 6607 9091 6613
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 10318 6604 10324 6656
rect 10376 6644 10382 6656
rect 12069 6647 12127 6653
rect 12069 6644 12081 6647
rect 10376 6616 12081 6644
rect 10376 6604 10382 6616
rect 12069 6613 12081 6616
rect 12115 6613 12127 6647
rect 13170 6644 13176 6656
rect 13131 6616 13176 6644
rect 12069 6607 12127 6613
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 5074 6400 5080 6452
rect 5132 6440 5138 6452
rect 8018 6440 8024 6452
rect 5132 6412 8024 6440
rect 5132 6400 5138 6412
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 9582 6440 9588 6452
rect 8168 6412 9588 6440
rect 8168 6400 8174 6412
rect 9582 6400 9588 6412
rect 9640 6440 9646 6452
rect 12434 6440 12440 6452
rect 9640 6412 10364 6440
rect 12395 6412 12440 6440
rect 9640 6400 9646 6412
rect 5353 6375 5411 6381
rect 5353 6341 5365 6375
rect 5399 6341 5411 6375
rect 5353 6335 5411 6341
rect 9401 6375 9459 6381
rect 9401 6341 9413 6375
rect 9447 6372 9459 6375
rect 9858 6372 9864 6384
rect 9447 6344 9864 6372
rect 9447 6341 9459 6344
rect 9401 6335 9459 6341
rect 1946 6304 1952 6316
rect 1859 6276 1952 6304
rect 1946 6264 1952 6276
rect 2004 6304 2010 6316
rect 2590 6304 2596 6316
rect 2004 6276 2596 6304
rect 2004 6264 2010 6276
rect 2590 6264 2596 6276
rect 2648 6264 2654 6316
rect 4062 6304 4068 6316
rect 4023 6276 4068 6304
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6304 4767 6307
rect 4982 6304 4988 6316
rect 4755 6276 4988 6304
rect 4755 6273 4767 6276
rect 4709 6267 4767 6273
rect 4982 6264 4988 6276
rect 5040 6264 5046 6316
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6304 5227 6307
rect 5258 6304 5264 6316
rect 5215 6276 5264 6304
rect 5215 6273 5227 6276
rect 5169 6267 5227 6273
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 5368 6302 5396 6335
rect 9858 6332 9864 6344
rect 9916 6372 9922 6384
rect 10226 6372 10232 6384
rect 9916 6344 10232 6372
rect 9916 6332 9922 6344
rect 10226 6332 10232 6344
rect 10284 6332 10290 6384
rect 10336 6372 10364 6412
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 13265 6375 13323 6381
rect 13265 6372 13277 6375
rect 10336 6344 13277 6372
rect 13265 6341 13277 6344
rect 13311 6341 13323 6375
rect 46382 6372 46388 6384
rect 13265 6335 13323 6341
rect 45204 6344 46388 6372
rect 5368 6274 5488 6302
rect 3602 6168 3608 6180
rect 2792 6140 3608 6168
rect 1670 6060 1676 6112
rect 1728 6100 1734 6112
rect 2041 6103 2099 6109
rect 2041 6100 2053 6103
rect 1728 6072 2053 6100
rect 1728 6060 1734 6072
rect 2041 6069 2053 6072
rect 2087 6069 2099 6103
rect 2041 6063 2099 6069
rect 2685 6103 2743 6109
rect 2685 6069 2697 6103
rect 2731 6100 2743 6103
rect 2792 6100 2820 6140
rect 3602 6128 3608 6140
rect 3660 6128 3666 6180
rect 4525 6171 4583 6177
rect 4525 6137 4537 6171
rect 4571 6168 4583 6171
rect 4982 6168 4988 6180
rect 4571 6140 4988 6168
rect 4571 6137 4583 6140
rect 4525 6131 4583 6137
rect 4982 6128 4988 6140
rect 5040 6168 5046 6180
rect 5460 6168 5488 6274
rect 5718 6264 5724 6316
rect 5776 6304 5782 6316
rect 6362 6304 6368 6316
rect 5776 6276 6368 6304
rect 5776 6264 5782 6276
rect 6362 6264 6368 6276
rect 6420 6264 6426 6316
rect 7742 6264 7748 6316
rect 7800 6264 7806 6316
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6304 8631 6307
rect 8938 6304 8944 6316
rect 8619 6276 8944 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 9490 6264 9496 6316
rect 9548 6304 9554 6316
rect 9585 6307 9643 6313
rect 9585 6304 9597 6307
rect 9548 6276 9597 6304
rect 9548 6264 9554 6276
rect 9585 6273 9597 6276
rect 9631 6273 9643 6307
rect 9585 6267 9643 6273
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 10318 6304 10324 6316
rect 9732 6276 9777 6304
rect 10279 6276 10324 6304
rect 9732 6264 9738 6276
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 12342 6304 12348 6316
rect 12303 6276 12348 6304
rect 12342 6264 12348 6276
rect 12400 6304 12406 6316
rect 13081 6307 13139 6313
rect 13081 6304 13093 6307
rect 12400 6276 13093 6304
rect 12400 6264 12406 6276
rect 13081 6273 13093 6276
rect 13127 6273 13139 6307
rect 13081 6267 13139 6273
rect 13725 6307 13783 6313
rect 13725 6273 13737 6307
rect 13771 6304 13783 6307
rect 14366 6304 14372 6316
rect 13771 6276 14372 6304
rect 13771 6273 13783 6276
rect 13725 6267 13783 6273
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 45204 6313 45232 6344
rect 46382 6332 46388 6344
rect 46440 6332 46446 6384
rect 45189 6307 45247 6313
rect 45189 6273 45201 6307
rect 45235 6273 45247 6307
rect 45189 6267 45247 6273
rect 6638 6236 6644 6248
rect 6599 6208 6644 6236
rect 6638 6196 6644 6208
rect 6696 6196 6702 6248
rect 6730 6196 6736 6248
rect 6788 6236 6794 6248
rect 6788 6208 8800 6236
rect 6788 6196 6794 6208
rect 5040 6140 5488 6168
rect 5040 6128 5046 6140
rect 3418 6100 3424 6112
rect 2731 6072 2820 6100
rect 3379 6072 3424 6100
rect 2731 6069 2743 6072
rect 2685 6063 2743 6069
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 3881 6103 3939 6109
rect 3881 6069 3893 6103
rect 3927 6100 3939 6103
rect 3970 6100 3976 6112
rect 3927 6072 3976 6100
rect 3927 6069 3939 6072
rect 3881 6063 3939 6069
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 4890 6060 4896 6112
rect 4948 6100 4954 6112
rect 5537 6103 5595 6109
rect 5537 6100 5549 6103
rect 4948 6072 5549 6100
rect 4948 6060 4954 6072
rect 5537 6069 5549 6072
rect 5583 6069 5595 6103
rect 5537 6063 5595 6069
rect 7098 6060 7104 6112
rect 7156 6100 7162 6112
rect 8113 6103 8171 6109
rect 8113 6100 8125 6103
rect 7156 6072 8125 6100
rect 7156 6060 7162 6072
rect 8113 6069 8125 6072
rect 8159 6069 8171 6103
rect 8662 6100 8668 6112
rect 8623 6072 8668 6100
rect 8113 6063 8171 6069
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 8772 6100 8800 6208
rect 9766 6196 9772 6248
rect 9824 6236 9830 6248
rect 10413 6239 10471 6245
rect 10413 6236 10425 6239
rect 9824 6208 10425 6236
rect 9824 6196 9830 6208
rect 10413 6205 10425 6208
rect 10459 6205 10471 6239
rect 10413 6199 10471 6205
rect 9398 6168 9404 6180
rect 9359 6140 9404 6168
rect 9398 6128 9404 6140
rect 9456 6128 9462 6180
rect 10428 6168 10456 6199
rect 10594 6196 10600 6248
rect 10652 6236 10658 6248
rect 10689 6239 10747 6245
rect 10689 6236 10701 6239
rect 10652 6208 10701 6236
rect 10652 6196 10658 6208
rect 10689 6205 10701 6208
rect 10735 6205 10747 6239
rect 45370 6236 45376 6248
rect 45331 6208 45376 6236
rect 10689 6199 10747 6205
rect 45370 6196 45376 6208
rect 45428 6196 45434 6248
rect 47029 6239 47087 6245
rect 47029 6205 47041 6239
rect 47075 6236 47087 6239
rect 48406 6236 48412 6248
rect 47075 6208 48412 6236
rect 47075 6205 47087 6208
rect 47029 6199 47087 6205
rect 48406 6196 48412 6208
rect 48464 6196 48470 6248
rect 11790 6168 11796 6180
rect 10428 6140 11796 6168
rect 11790 6128 11796 6140
rect 11848 6128 11854 6180
rect 13446 6128 13452 6180
rect 13504 6168 13510 6180
rect 14461 6171 14519 6177
rect 14461 6168 14473 6171
rect 13504 6140 14473 6168
rect 13504 6128 13510 6140
rect 14461 6137 14473 6140
rect 14507 6137 14519 6171
rect 14461 6131 14519 6137
rect 12434 6100 12440 6112
rect 8772 6072 12440 6100
rect 12434 6060 12440 6072
rect 12492 6060 12498 6112
rect 13814 6100 13820 6112
rect 13775 6072 13820 6100
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 46290 6060 46296 6112
rect 46348 6100 46354 6112
rect 47765 6103 47823 6109
rect 47765 6100 47777 6103
rect 46348 6072 47777 6100
rect 46348 6060 46354 6072
rect 47765 6069 47777 6072
rect 47811 6069 47823 6103
rect 47765 6063 47823 6069
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 3881 5899 3939 5905
rect 3881 5865 3893 5899
rect 3927 5896 3939 5899
rect 6270 5896 6276 5908
rect 3927 5868 6276 5896
rect 3927 5865 3939 5868
rect 3881 5859 3939 5865
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 10226 5856 10232 5908
rect 10284 5896 10290 5908
rect 11609 5899 11667 5905
rect 11609 5896 11621 5899
rect 10284 5868 11621 5896
rect 10284 5856 10290 5868
rect 11609 5865 11621 5868
rect 11655 5865 11667 5899
rect 11790 5896 11796 5908
rect 11751 5868 11796 5896
rect 11609 5859 11667 5865
rect 11790 5856 11796 5868
rect 11848 5856 11854 5908
rect 12434 5896 12440 5908
rect 12395 5868 12440 5896
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 8386 5788 8392 5840
rect 8444 5828 8450 5840
rect 9493 5831 9551 5837
rect 9493 5828 9505 5831
rect 8444 5800 9505 5828
rect 8444 5788 8450 5800
rect 9493 5797 9505 5800
rect 9539 5797 9551 5831
rect 12342 5828 12348 5840
rect 12255 5800 12348 5828
rect 9493 5791 9551 5797
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5760 2007 5763
rect 3234 5760 3240 5772
rect 1995 5732 3240 5760
rect 1995 5729 2007 5732
rect 1949 5723 2007 5729
rect 3234 5720 3240 5732
rect 3292 5720 3298 5772
rect 7282 5760 7288 5772
rect 5828 5732 7288 5760
rect 2409 5695 2467 5701
rect 2409 5661 2421 5695
rect 2455 5692 2467 5695
rect 3053 5695 3111 5701
rect 3053 5692 3065 5695
rect 2455 5664 3065 5692
rect 2455 5661 2467 5664
rect 2409 5655 2467 5661
rect 3053 5661 3065 5664
rect 3099 5692 3111 5695
rect 3326 5692 3332 5704
rect 3099 5664 3332 5692
rect 3099 5661 3111 5664
rect 3053 5655 3111 5661
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 3694 5652 3700 5704
rect 3752 5692 3758 5704
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 3752 5664 3801 5692
rect 3752 5652 3758 5664
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 4430 5692 4436 5704
rect 4391 5664 4436 5692
rect 3789 5655 3847 5661
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 5828 5678 5856 5732
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 7558 5720 7564 5772
rect 7616 5760 7622 5772
rect 9033 5763 9091 5769
rect 9033 5760 9045 5763
rect 7616 5732 9045 5760
rect 7616 5720 7622 5732
rect 9033 5729 9045 5732
rect 9079 5760 9091 5763
rect 9674 5760 9680 5772
rect 9079 5732 9680 5760
rect 9079 5729 9091 5732
rect 9033 5723 9091 5729
rect 9674 5720 9680 5732
rect 9732 5760 9738 5772
rect 10502 5760 10508 5772
rect 9732 5732 10508 5760
rect 9732 5720 9738 5732
rect 10502 5720 10508 5732
rect 10560 5720 10566 5772
rect 10686 5760 10692 5772
rect 10647 5732 10692 5760
rect 10686 5720 10692 5732
rect 10744 5720 10750 5772
rect 10965 5763 11023 5769
rect 10965 5729 10977 5763
rect 11011 5760 11023 5763
rect 11790 5760 11796 5772
rect 11011 5732 11796 5760
rect 11011 5729 11023 5732
rect 10965 5723 11023 5729
rect 11790 5720 11796 5732
rect 11848 5720 11854 5772
rect 6362 5652 6368 5704
rect 6420 5692 6426 5704
rect 6641 5695 6699 5701
rect 6641 5692 6653 5695
rect 6420 5664 6653 5692
rect 6420 5652 6426 5664
rect 6641 5661 6653 5664
rect 6687 5661 6699 5695
rect 8662 5692 8668 5704
rect 8050 5664 8668 5692
rect 6641 5655 6699 5661
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5692 9183 5695
rect 9490 5692 9496 5704
rect 9171 5664 9496 5692
rect 9171 5661 9183 5664
rect 9125 5655 9183 5661
rect 9490 5652 9496 5664
rect 9548 5652 9554 5704
rect 9582 5652 9588 5704
rect 9640 5692 9646 5704
rect 12268 5701 12296 5800
rect 12342 5788 12348 5800
rect 12400 5828 12406 5840
rect 13906 5828 13912 5840
rect 12400 5800 13912 5828
rect 12400 5788 12406 5800
rect 13906 5788 13912 5800
rect 13964 5788 13970 5840
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 15013 5763 15071 5769
rect 15013 5760 15025 5763
rect 12492 5732 15025 5760
rect 12492 5720 12498 5732
rect 15013 5729 15025 5732
rect 15059 5729 15071 5763
rect 15013 5723 15071 5729
rect 31021 5763 31079 5769
rect 31021 5729 31033 5763
rect 31067 5760 31079 5763
rect 31846 5760 31852 5772
rect 31067 5732 31852 5760
rect 31067 5729 31079 5732
rect 31021 5723 31079 5729
rect 31846 5720 31852 5732
rect 31904 5720 31910 5772
rect 44453 5763 44511 5769
rect 44453 5729 44465 5763
rect 44499 5760 44511 5763
rect 45830 5760 45836 5772
rect 44499 5732 45836 5760
rect 44499 5729 44511 5732
rect 44453 5723 44511 5729
rect 45830 5720 45836 5732
rect 45888 5720 45894 5772
rect 46290 5760 46296 5772
rect 46251 5732 46296 5760
rect 46290 5720 46296 5732
rect 46348 5720 46354 5772
rect 47118 5760 47124 5772
rect 47079 5732 47124 5760
rect 47118 5720 47124 5732
rect 47176 5720 47182 5772
rect 10597 5695 10655 5701
rect 10597 5692 10609 5695
rect 9640 5664 10609 5692
rect 9640 5652 9646 5664
rect 10597 5661 10609 5664
rect 10643 5661 10655 5695
rect 10597 5655 10655 5661
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5661 12311 5695
rect 12253 5655 12311 5661
rect 13357 5695 13415 5701
rect 13357 5661 13369 5695
rect 13403 5692 13415 5695
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 13403 5664 14289 5692
rect 13403 5661 13415 5664
rect 13357 5655 13415 5661
rect 14277 5661 14289 5664
rect 14323 5692 14335 5695
rect 14366 5692 14372 5704
rect 14323 5664 14372 5692
rect 14323 5661 14335 5664
rect 14277 5655 14335 5661
rect 14366 5652 14372 5664
rect 14424 5692 14430 5704
rect 14918 5692 14924 5704
rect 14424 5664 14924 5692
rect 14424 5652 14430 5664
rect 14918 5652 14924 5664
rect 14976 5652 14982 5704
rect 31665 5695 31723 5701
rect 31665 5661 31677 5695
rect 31711 5692 31723 5695
rect 31938 5692 31944 5704
rect 31711 5664 31944 5692
rect 31711 5661 31723 5664
rect 31665 5655 31723 5661
rect 31938 5652 31944 5664
rect 31996 5652 32002 5704
rect 32122 5652 32128 5704
rect 32180 5692 32186 5704
rect 32309 5695 32367 5701
rect 32309 5692 32321 5695
rect 32180 5664 32321 5692
rect 32180 5652 32186 5664
rect 32309 5661 32321 5664
rect 32355 5661 32367 5695
rect 36354 5692 36360 5704
rect 36315 5664 36360 5692
rect 32309 5655 32367 5661
rect 36354 5652 36360 5664
rect 36412 5652 36418 5704
rect 37001 5695 37059 5701
rect 37001 5661 37013 5695
rect 37047 5692 37059 5695
rect 37274 5692 37280 5704
rect 37047 5664 37280 5692
rect 37047 5661 37059 5664
rect 37001 5655 37059 5661
rect 37274 5652 37280 5664
rect 37332 5652 37338 5704
rect 38381 5695 38439 5701
rect 38381 5661 38393 5695
rect 38427 5692 38439 5695
rect 39574 5692 39580 5704
rect 38427 5664 39580 5692
rect 38427 5661 38439 5664
rect 38381 5655 38439 5661
rect 39574 5652 39580 5664
rect 39632 5652 39638 5704
rect 40126 5652 40132 5704
rect 40184 5692 40190 5704
rect 40221 5695 40279 5701
rect 40221 5692 40233 5695
rect 40184 5664 40233 5692
rect 40184 5652 40190 5664
rect 40221 5661 40233 5664
rect 40267 5661 40279 5695
rect 41598 5692 41604 5704
rect 41559 5664 41604 5692
rect 40221 5655 40279 5661
rect 41598 5652 41604 5664
rect 41656 5652 41662 5704
rect 43349 5695 43407 5701
rect 43349 5661 43361 5695
rect 43395 5692 43407 5695
rect 45002 5692 45008 5704
rect 43395 5664 45008 5692
rect 43395 5661 43407 5664
rect 43349 5655 43407 5661
rect 45002 5652 45008 5664
rect 45060 5652 45066 5704
rect 45646 5692 45652 5704
rect 45607 5664 45652 5692
rect 45646 5652 45652 5664
rect 45704 5652 45710 5704
rect 3145 5627 3203 5633
rect 3145 5593 3157 5627
rect 3191 5624 3203 5627
rect 4246 5624 4252 5636
rect 3191 5596 4252 5624
rect 3191 5593 3203 5596
rect 3145 5587 3203 5593
rect 4246 5584 4252 5596
rect 4304 5584 4310 5636
rect 4614 5584 4620 5636
rect 4672 5624 4678 5636
rect 4709 5627 4767 5633
rect 4709 5624 4721 5627
rect 4672 5596 4721 5624
rect 4672 5584 4678 5596
rect 4709 5593 4721 5596
rect 4755 5593 4767 5627
rect 6917 5627 6975 5633
rect 6917 5624 6929 5627
rect 4709 5587 4767 5593
rect 6012 5596 6929 5624
rect 2501 5559 2559 5565
rect 2501 5525 2513 5559
rect 2547 5556 2559 5559
rect 3786 5556 3792 5568
rect 2547 5528 3792 5556
rect 2547 5525 2559 5528
rect 2501 5519 2559 5525
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 4154 5516 4160 5568
rect 4212 5556 4218 5568
rect 6012 5556 6040 5596
rect 6917 5593 6929 5596
rect 6963 5593 6975 5627
rect 9508 5624 9536 5652
rect 11425 5627 11483 5633
rect 11425 5624 11437 5627
rect 9508 5596 11437 5624
rect 6917 5587 6975 5593
rect 11425 5593 11437 5596
rect 11471 5593 11483 5627
rect 11425 5587 11483 5593
rect 12158 5584 12164 5636
rect 12216 5624 12222 5636
rect 13449 5627 13507 5633
rect 13449 5624 13461 5627
rect 12216 5596 13461 5624
rect 12216 5584 12222 5596
rect 13449 5593 13461 5596
rect 13495 5593 13507 5627
rect 13449 5587 13507 5593
rect 45741 5627 45799 5633
rect 45741 5593 45753 5627
rect 45787 5624 45799 5627
rect 46477 5627 46535 5633
rect 46477 5624 46489 5627
rect 45787 5596 46489 5624
rect 45787 5593 45799 5596
rect 45741 5587 45799 5593
rect 46477 5593 46489 5596
rect 46523 5593 46535 5627
rect 46477 5587 46535 5593
rect 6178 5556 6184 5568
rect 4212 5528 6040 5556
rect 6139 5528 6184 5556
rect 4212 5516 4218 5528
rect 6178 5516 6184 5528
rect 6236 5556 6242 5568
rect 6822 5556 6828 5568
rect 6236 5528 6828 5556
rect 6236 5516 6242 5528
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 7190 5516 7196 5568
rect 7248 5556 7254 5568
rect 8389 5559 8447 5565
rect 8389 5556 8401 5559
rect 7248 5528 8401 5556
rect 7248 5516 7254 5528
rect 8389 5525 8401 5528
rect 8435 5525 8447 5559
rect 8389 5519 8447 5525
rect 10502 5516 10508 5568
rect 10560 5556 10566 5568
rect 11625 5559 11683 5565
rect 11625 5556 11637 5559
rect 10560 5528 11637 5556
rect 10560 5516 10566 5528
rect 11625 5525 11637 5528
rect 11671 5525 11683 5559
rect 11625 5519 11683 5525
rect 14369 5559 14427 5565
rect 14369 5525 14381 5559
rect 14415 5556 14427 5559
rect 14458 5556 14464 5568
rect 14415 5528 14464 5556
rect 14415 5525 14427 5528
rect 14369 5519 14427 5525
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 43441 5559 43499 5565
rect 43441 5525 43453 5559
rect 43487 5556 43499 5559
rect 44910 5556 44916 5568
rect 43487 5528 44916 5556
rect 43487 5525 43499 5528
rect 43441 5519 43499 5525
rect 44910 5516 44916 5528
rect 44968 5516 44974 5568
rect 45097 5559 45155 5565
rect 45097 5525 45109 5559
rect 45143 5556 45155 5559
rect 45186 5556 45192 5568
rect 45143 5528 45192 5556
rect 45143 5525 45155 5528
rect 45097 5519 45155 5525
rect 45186 5516 45192 5528
rect 45244 5516 45250 5568
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 3605 5355 3663 5361
rect 3605 5321 3617 5355
rect 3651 5352 3663 5355
rect 4154 5352 4160 5364
rect 3651 5324 4160 5352
rect 3651 5321 3663 5324
rect 3605 5315 3663 5321
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 4801 5355 4859 5361
rect 4801 5321 4813 5355
rect 4847 5352 4859 5355
rect 6638 5352 6644 5364
rect 4847 5324 6644 5352
rect 4847 5321 4859 5324
rect 4801 5315 4859 5321
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 6822 5312 6828 5364
rect 6880 5352 6886 5364
rect 7009 5355 7067 5361
rect 7009 5352 7021 5355
rect 6880 5324 7021 5352
rect 6880 5312 6886 5324
rect 7009 5321 7021 5324
rect 7055 5321 7067 5355
rect 7190 5352 7196 5364
rect 7151 5324 7196 5352
rect 7009 5315 7067 5321
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 7377 5355 7435 5361
rect 7377 5321 7389 5355
rect 7423 5352 7435 5355
rect 7558 5352 7564 5364
rect 7423 5324 7564 5352
rect 7423 5321 7435 5324
rect 7377 5315 7435 5321
rect 7558 5312 7564 5324
rect 7616 5312 7622 5364
rect 10318 5312 10324 5364
rect 10376 5352 10382 5364
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 10376 5324 10425 5352
rect 10376 5312 10382 5324
rect 10413 5321 10425 5324
rect 10459 5321 10471 5355
rect 10413 5315 10471 5321
rect 10502 5312 10508 5364
rect 10560 5352 10566 5364
rect 10686 5352 10692 5364
rect 10560 5324 10605 5352
rect 10647 5324 10692 5352
rect 10560 5312 10566 5324
rect 10686 5312 10692 5324
rect 10744 5312 10750 5364
rect 13265 5355 13323 5361
rect 13265 5352 13277 5355
rect 10796 5324 13277 5352
rect 2409 5287 2467 5293
rect 2409 5253 2421 5287
rect 2455 5284 2467 5287
rect 2590 5284 2596 5296
rect 2455 5256 2596 5284
rect 2455 5253 2467 5256
rect 2409 5247 2467 5253
rect 2590 5244 2596 5256
rect 2648 5244 2654 5296
rect 5074 5284 5080 5296
rect 3804 5256 5080 5284
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5216 2283 5219
rect 2314 5216 2320 5228
rect 2271 5188 2320 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 2682 5176 2688 5228
rect 2740 5216 2746 5228
rect 2961 5219 3019 5225
rect 2961 5216 2973 5219
rect 2740 5188 2973 5216
rect 2740 5176 2746 5188
rect 2961 5185 2973 5188
rect 3007 5216 3019 5219
rect 3694 5216 3700 5228
rect 3007 5188 3700 5216
rect 3007 5185 3019 5188
rect 2961 5179 3019 5185
rect 3694 5176 3700 5188
rect 3752 5176 3758 5228
rect 3804 5225 3832 5256
rect 5074 5244 5080 5256
rect 5132 5244 5138 5296
rect 7098 5284 7104 5296
rect 5460 5256 7104 5284
rect 5460 5225 5488 5256
rect 7098 5244 7104 5256
rect 7156 5244 7162 5296
rect 8113 5287 8171 5293
rect 8113 5253 8125 5287
rect 8159 5284 8171 5287
rect 8386 5284 8392 5296
rect 8159 5256 8392 5284
rect 8159 5253 8171 5256
rect 8113 5247 8171 5253
rect 8386 5244 8392 5256
rect 8444 5244 8450 5296
rect 9122 5244 9128 5296
rect 9180 5244 9186 5296
rect 9582 5244 9588 5296
rect 9640 5284 9646 5296
rect 10796 5284 10824 5324
rect 13265 5321 13277 5324
rect 13311 5321 13323 5355
rect 13265 5315 13323 5321
rect 11790 5284 11796 5296
rect 9640 5256 10824 5284
rect 11751 5256 11796 5284
rect 9640 5244 9646 5256
rect 11790 5244 11796 5256
rect 11848 5244 11854 5296
rect 13170 5284 13176 5296
rect 13018 5256 13176 5284
rect 13170 5244 13176 5256
rect 13228 5244 13234 5296
rect 45462 5284 45468 5296
rect 45204 5256 45468 5284
rect 3789 5219 3847 5225
rect 3789 5185 3801 5219
rect 3835 5185 3847 5219
rect 3789 5179 3847 5185
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5216 4491 5219
rect 5445 5219 5503 5225
rect 5445 5216 5457 5219
rect 4479 5188 5457 5216
rect 4479 5185 4491 5188
rect 4433 5179 4491 5185
rect 5445 5185 5457 5188
rect 5491 5185 5503 5219
rect 5626 5216 5632 5228
rect 5587 5188 5632 5216
rect 5445 5179 5503 5185
rect 5626 5176 5632 5188
rect 5684 5216 5690 5228
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 5684 5188 6837 5216
rect 5684 5176 5690 5188
rect 6825 5185 6837 5188
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 10226 5176 10232 5228
rect 10284 5216 10290 5228
rect 10321 5219 10379 5225
rect 10321 5216 10333 5219
rect 10284 5188 10333 5216
rect 10284 5176 10290 5188
rect 10321 5185 10333 5188
rect 10367 5185 10379 5219
rect 10321 5179 10379 5185
rect 16482 5176 16488 5228
rect 16540 5216 16546 5228
rect 16669 5219 16727 5225
rect 16669 5216 16681 5219
rect 16540 5188 16681 5216
rect 16540 5176 16546 5188
rect 16669 5185 16681 5188
rect 16715 5216 16727 5219
rect 17313 5219 17371 5225
rect 17313 5216 17325 5219
rect 16715 5188 17325 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 17313 5185 17325 5188
rect 17359 5216 17371 5219
rect 18325 5219 18383 5225
rect 18325 5216 18337 5219
rect 17359 5188 18337 5216
rect 17359 5185 17371 5188
rect 17313 5179 17371 5185
rect 18325 5185 18337 5188
rect 18371 5185 18383 5219
rect 18325 5179 18383 5185
rect 18414 5176 18420 5228
rect 18472 5216 18478 5228
rect 20257 5219 20315 5225
rect 20257 5216 20269 5219
rect 18472 5188 20269 5216
rect 18472 5176 18478 5188
rect 20257 5185 20269 5188
rect 20303 5216 20315 5219
rect 21082 5216 21088 5228
rect 20303 5188 21088 5216
rect 20303 5185 20315 5188
rect 20257 5179 20315 5185
rect 21082 5176 21088 5188
rect 21140 5216 21146 5228
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 21140 5188 21833 5216
rect 21140 5176 21146 5188
rect 21821 5185 21833 5188
rect 21867 5185 21879 5219
rect 21821 5179 21879 5185
rect 28353 5219 28411 5225
rect 28353 5185 28365 5219
rect 28399 5216 28411 5219
rect 28534 5216 28540 5228
rect 28399 5188 28540 5216
rect 28399 5185 28411 5188
rect 28353 5179 28411 5185
rect 28534 5176 28540 5188
rect 28592 5216 28598 5228
rect 28997 5219 29055 5225
rect 28997 5216 29009 5219
rect 28592 5188 29009 5216
rect 28592 5176 28598 5188
rect 28997 5185 29009 5188
rect 29043 5185 29055 5219
rect 28997 5179 29055 5185
rect 30469 5219 30527 5225
rect 30469 5185 30481 5219
rect 30515 5216 30527 5219
rect 31113 5219 31171 5225
rect 31113 5216 31125 5219
rect 30515 5188 31125 5216
rect 30515 5185 30527 5188
rect 30469 5179 30527 5185
rect 31113 5185 31125 5188
rect 31159 5216 31171 5219
rect 31662 5216 31668 5228
rect 31159 5188 31668 5216
rect 31159 5185 31171 5188
rect 31113 5179 31171 5185
rect 31662 5176 31668 5188
rect 31720 5216 31726 5228
rect 32125 5219 32183 5225
rect 32125 5216 32137 5219
rect 31720 5188 32137 5216
rect 31720 5176 31726 5188
rect 32125 5185 32137 5188
rect 32171 5216 32183 5219
rect 32769 5219 32827 5225
rect 32769 5216 32781 5219
rect 32171 5188 32781 5216
rect 32171 5185 32183 5188
rect 32125 5179 32183 5185
rect 32769 5185 32781 5188
rect 32815 5185 32827 5219
rect 33410 5216 33416 5228
rect 33371 5188 33416 5216
rect 32769 5179 32827 5185
rect 33410 5176 33416 5188
rect 33468 5216 33474 5228
rect 34057 5219 34115 5225
rect 34057 5216 34069 5219
rect 33468 5188 34069 5216
rect 33468 5176 33474 5188
rect 34057 5185 34069 5188
rect 34103 5216 34115 5219
rect 35345 5219 35403 5225
rect 35345 5216 35357 5219
rect 34103 5188 35357 5216
rect 34103 5185 34115 5188
rect 34057 5179 34115 5185
rect 35345 5185 35357 5188
rect 35391 5216 35403 5219
rect 35434 5216 35440 5228
rect 35391 5188 35440 5216
rect 35391 5185 35403 5188
rect 35345 5179 35403 5185
rect 35434 5176 35440 5188
rect 35492 5176 35498 5228
rect 37277 5219 37335 5225
rect 37277 5185 37289 5219
rect 37323 5216 37335 5219
rect 37918 5216 37924 5228
rect 37323 5188 37924 5216
rect 37323 5185 37335 5188
rect 37277 5179 37335 5185
rect 37918 5176 37924 5188
rect 37976 5216 37982 5228
rect 38565 5219 38623 5225
rect 38565 5216 38577 5219
rect 37976 5188 38577 5216
rect 37976 5176 37982 5188
rect 38565 5185 38577 5188
rect 38611 5185 38623 5219
rect 38565 5179 38623 5185
rect 40497 5219 40555 5225
rect 40497 5185 40509 5219
rect 40543 5216 40555 5219
rect 41141 5219 41199 5225
rect 41141 5216 41153 5219
rect 40543 5188 41153 5216
rect 40543 5185 40555 5188
rect 40497 5179 40555 5185
rect 41141 5185 41153 5188
rect 41187 5216 41199 5219
rect 42426 5216 42432 5228
rect 41187 5188 42432 5216
rect 41187 5185 41199 5188
rect 41141 5179 41199 5185
rect 42426 5176 42432 5188
rect 42484 5176 42490 5228
rect 43717 5219 43775 5225
rect 43717 5185 43729 5219
rect 43763 5216 43775 5219
rect 44361 5219 44419 5225
rect 44361 5216 44373 5219
rect 43763 5188 44373 5216
rect 43763 5185 43775 5188
rect 43717 5179 43775 5185
rect 44361 5185 44373 5188
rect 44407 5216 44419 5219
rect 45002 5216 45008 5228
rect 44407 5188 45008 5216
rect 44407 5185 44419 5188
rect 44361 5179 44419 5185
rect 45002 5176 45008 5188
rect 45060 5176 45066 5228
rect 45204 5225 45232 5256
rect 45462 5244 45468 5256
rect 45520 5244 45526 5296
rect 45189 5219 45247 5225
rect 45189 5185 45201 5219
rect 45235 5185 45247 5219
rect 47578 5216 47584 5228
rect 45189 5179 45247 5185
rect 46768 5188 47584 5216
rect 2866 5108 2872 5160
rect 2924 5148 2930 5160
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 2924 5120 4353 5148
rect 2924 5108 2930 5120
rect 4341 5117 4353 5120
rect 4387 5117 4399 5151
rect 5534 5148 5540 5160
rect 5495 5120 5540 5148
rect 4341 5111 4399 5117
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 6546 5148 6552 5160
rect 5767 5120 6552 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 6546 5108 6552 5120
rect 6604 5148 6610 5160
rect 7190 5148 7196 5160
rect 6604 5120 7196 5148
rect 6604 5108 6610 5120
rect 7190 5108 7196 5120
rect 7248 5108 7254 5160
rect 7837 5151 7895 5157
rect 7837 5117 7849 5151
rect 7883 5148 7895 5151
rect 8478 5148 8484 5160
rect 7883 5120 8484 5148
rect 7883 5117 7895 5120
rect 7837 5111 7895 5117
rect 8478 5108 8484 5120
rect 8536 5148 8542 5160
rect 11517 5151 11575 5157
rect 11517 5148 11529 5151
rect 8536 5120 11529 5148
rect 8536 5108 8542 5120
rect 11517 5117 11529 5120
rect 11563 5117 11575 5151
rect 45370 5148 45376 5160
rect 45331 5120 45376 5148
rect 11517 5111 11575 5117
rect 45370 5108 45376 5120
rect 45428 5108 45434 5160
rect 45646 5108 45652 5160
rect 45704 5148 45710 5160
rect 46768 5148 46796 5188
rect 47578 5176 47584 5188
rect 47636 5176 47642 5228
rect 45704 5120 46796 5148
rect 47029 5151 47087 5157
rect 45704 5108 45710 5120
rect 47029 5117 47041 5151
rect 47075 5148 47087 5151
rect 47670 5148 47676 5160
rect 47075 5120 47676 5148
rect 47075 5117 47087 5120
rect 47029 5111 47087 5117
rect 47670 5108 47676 5120
rect 47728 5108 47734 5160
rect 1673 5083 1731 5089
rect 1673 5049 1685 5083
rect 1719 5080 1731 5083
rect 3970 5080 3976 5092
rect 1719 5052 3976 5080
rect 1719 5049 1731 5052
rect 1673 5043 1731 5049
rect 3970 5040 3976 5052
rect 4028 5040 4034 5092
rect 5261 5083 5319 5089
rect 5261 5049 5273 5083
rect 5307 5080 5319 5083
rect 5810 5080 5816 5092
rect 5307 5052 5816 5080
rect 5307 5049 5319 5052
rect 5261 5043 5319 5049
rect 5810 5040 5816 5052
rect 5868 5040 5874 5092
rect 10137 5083 10195 5089
rect 10137 5049 10149 5083
rect 10183 5049 10195 5083
rect 10137 5043 10195 5049
rect 3050 5012 3056 5024
rect 3011 4984 3056 5012
rect 3050 4972 3056 4984
rect 3108 4972 3114 5024
rect 9490 4972 9496 5024
rect 9548 5012 9554 5024
rect 9585 5015 9643 5021
rect 9585 5012 9597 5015
rect 9548 4984 9597 5012
rect 9548 4972 9554 4984
rect 9585 4981 9597 4984
rect 9631 5012 9643 5015
rect 10152 5012 10180 5043
rect 14090 5040 14096 5092
rect 14148 5080 14154 5092
rect 15105 5083 15163 5089
rect 15105 5080 15117 5083
rect 14148 5052 15117 5080
rect 14148 5040 14154 5052
rect 15105 5049 15117 5052
rect 15151 5049 15163 5083
rect 15105 5043 15163 5049
rect 30561 5083 30619 5089
rect 30561 5049 30573 5083
rect 30607 5080 30619 5083
rect 32398 5080 32404 5092
rect 30607 5052 32404 5080
rect 30607 5049 30619 5052
rect 30561 5043 30619 5049
rect 32398 5040 32404 5052
rect 32456 5040 32462 5092
rect 33505 5083 33563 5089
rect 33505 5049 33517 5083
rect 33551 5080 33563 5083
rect 34606 5080 34612 5092
rect 33551 5052 34612 5080
rect 33551 5049 33563 5052
rect 33505 5043 33563 5049
rect 34606 5040 34612 5052
rect 34664 5040 34670 5092
rect 36173 5083 36231 5089
rect 36173 5049 36185 5083
rect 36219 5080 36231 5083
rect 37642 5080 37648 5092
rect 36219 5052 37648 5080
rect 36219 5049 36231 5052
rect 36173 5043 36231 5049
rect 37642 5040 37648 5052
rect 37700 5040 37706 5092
rect 14366 5012 14372 5024
rect 9631 4984 10180 5012
rect 14327 4984 14372 5012
rect 9631 4981 9643 4984
rect 9585 4975 9643 4981
rect 14366 4972 14372 4984
rect 14424 4972 14430 5024
rect 15194 4972 15200 5024
rect 15252 5012 15258 5024
rect 15749 5015 15807 5021
rect 15749 5012 15761 5015
rect 15252 4984 15761 5012
rect 15252 4972 15258 4984
rect 15749 4981 15761 4984
rect 15795 4981 15807 5015
rect 15749 4975 15807 4981
rect 15930 4972 15936 5024
rect 15988 5012 15994 5024
rect 16761 5015 16819 5021
rect 16761 5012 16773 5015
rect 15988 4984 16773 5012
rect 15988 4972 15994 4984
rect 16761 4981 16773 4984
rect 16807 4981 16819 5015
rect 17402 5012 17408 5024
rect 17363 4984 17408 5012
rect 16761 4975 16819 4981
rect 17402 4972 17408 4984
rect 17460 4972 17466 5024
rect 17954 4972 17960 5024
rect 18012 5012 18018 5024
rect 18417 5015 18475 5021
rect 18417 5012 18429 5015
rect 18012 4984 18429 5012
rect 18012 4972 18018 4984
rect 18417 4981 18429 4984
rect 18463 4981 18475 5015
rect 19150 5012 19156 5024
rect 19111 4984 19156 5012
rect 18417 4975 18475 4981
rect 19150 4972 19156 4984
rect 19208 4972 19214 5024
rect 19334 4972 19340 5024
rect 19392 5012 19398 5024
rect 19797 5015 19855 5021
rect 19797 5012 19809 5015
rect 19392 4984 19809 5012
rect 19392 4972 19398 4984
rect 19797 4981 19809 4984
rect 19843 4981 19855 5015
rect 20346 5012 20352 5024
rect 20307 4984 20352 5012
rect 19797 4975 19855 4981
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 20806 4972 20812 5024
rect 20864 5012 20870 5024
rect 21269 5015 21327 5021
rect 21269 5012 21281 5015
rect 20864 4984 21281 5012
rect 20864 4972 20870 4984
rect 21269 4981 21281 4984
rect 21315 4981 21327 5015
rect 21269 4975 21327 4981
rect 21450 4972 21456 5024
rect 21508 5012 21514 5024
rect 21913 5015 21971 5021
rect 21913 5012 21925 5015
rect 21508 4984 21925 5012
rect 21508 4972 21514 4984
rect 21913 4981 21925 4984
rect 21959 4981 21971 5015
rect 21913 4975 21971 4981
rect 22278 4972 22284 5024
rect 22336 5012 22342 5024
rect 23201 5015 23259 5021
rect 23201 5012 23213 5015
rect 22336 4984 23213 5012
rect 22336 4972 22342 4984
rect 23201 4981 23213 4984
rect 23247 4981 23259 5015
rect 23201 4975 23259 4981
rect 23842 4972 23848 5024
rect 23900 5012 23906 5024
rect 24121 5015 24179 5021
rect 24121 5012 24133 5015
rect 23900 4984 24133 5012
rect 23900 4972 23906 4984
rect 24121 4981 24133 4984
rect 24167 4981 24179 5015
rect 24121 4975 24179 4981
rect 24578 4972 24584 5024
rect 24636 5012 24642 5024
rect 24765 5015 24823 5021
rect 24765 5012 24777 5015
rect 24636 4984 24777 5012
rect 24636 4972 24642 4984
rect 24765 4981 24777 4984
rect 24811 4981 24823 5015
rect 28442 5012 28448 5024
rect 28403 4984 28448 5012
rect 24765 4975 24823 4981
rect 28442 4972 28448 4984
rect 28500 4972 28506 5024
rect 29086 5012 29092 5024
rect 29047 4984 29092 5012
rect 29086 4972 29092 4984
rect 29144 4972 29150 5024
rect 31205 5015 31263 5021
rect 31205 4981 31217 5015
rect 31251 5012 31263 5015
rect 32030 5012 32036 5024
rect 31251 4984 32036 5012
rect 31251 4981 31263 4984
rect 31205 4975 31263 4981
rect 32030 4972 32036 4984
rect 32088 4972 32094 5024
rect 32214 5012 32220 5024
rect 32175 4984 32220 5012
rect 32214 4972 32220 4984
rect 32272 4972 32278 5024
rect 32306 4972 32312 5024
rect 32364 5012 32370 5024
rect 32861 5015 32919 5021
rect 32861 5012 32873 5015
rect 32364 4984 32873 5012
rect 32364 4972 32370 4984
rect 32861 4981 32873 4984
rect 32907 4981 32919 5015
rect 32861 4975 32919 4981
rect 34149 5015 34207 5021
rect 34149 4981 34161 5015
rect 34195 5012 34207 5015
rect 34514 5012 34520 5024
rect 34195 4984 34520 5012
rect 34195 4981 34207 4984
rect 34149 4975 34207 4981
rect 34514 4972 34520 4984
rect 34572 4972 34578 5024
rect 34698 4972 34704 5024
rect 34756 5012 34762 5024
rect 34885 5015 34943 5021
rect 34885 5012 34897 5015
rect 34756 4984 34897 5012
rect 34756 4972 34762 4984
rect 34885 4981 34897 4984
rect 34931 4981 34943 5015
rect 34885 4975 34943 4981
rect 35342 4972 35348 5024
rect 35400 5012 35406 5024
rect 35437 5015 35495 5021
rect 35437 5012 35449 5015
rect 35400 4984 35449 5012
rect 35400 4972 35406 4984
rect 35437 4981 35449 4984
rect 35483 4981 35495 5015
rect 37366 5012 37372 5024
rect 37327 4984 37372 5012
rect 35437 4975 35495 4981
rect 37366 4972 37372 4984
rect 37424 4972 37430 5024
rect 37550 4972 37556 5024
rect 37608 5012 37614 5024
rect 38013 5015 38071 5021
rect 38013 5012 38025 5015
rect 37608 4984 38025 5012
rect 37608 4972 37614 4984
rect 38013 4981 38025 4984
rect 38059 4981 38071 5015
rect 38654 5012 38660 5024
rect 38615 4984 38660 5012
rect 38013 4975 38071 4981
rect 38654 4972 38660 4984
rect 38712 4972 38718 5024
rect 39390 5012 39396 5024
rect 39351 4984 39396 5012
rect 39390 4972 39396 4984
rect 39448 4972 39454 5024
rect 40037 5015 40095 5021
rect 40037 4981 40049 5015
rect 40083 5012 40095 5015
rect 40218 5012 40224 5024
rect 40083 4984 40224 5012
rect 40083 4981 40095 4984
rect 40037 4975 40095 4981
rect 40218 4972 40224 4984
rect 40276 4972 40282 5024
rect 40586 5012 40592 5024
rect 40547 4984 40592 5012
rect 40586 4972 40592 4984
rect 40644 4972 40650 5024
rect 41233 5015 41291 5021
rect 41233 4981 41245 5015
rect 41279 5012 41291 5015
rect 42058 5012 42064 5024
rect 41279 4984 42064 5012
rect 41279 4981 41291 4984
rect 41233 4975 41291 4981
rect 42058 4972 42064 4984
rect 42116 4972 42122 5024
rect 42521 5015 42579 5021
rect 42521 4981 42533 5015
rect 42567 5012 42579 5015
rect 42610 5012 42616 5024
rect 42567 4984 42616 5012
rect 42567 4981 42579 4984
rect 42521 4975 42579 4981
rect 42610 4972 42616 4984
rect 42668 4972 42674 5024
rect 43254 5012 43260 5024
rect 43215 4984 43260 5012
rect 43254 4972 43260 4984
rect 43312 4972 43318 5024
rect 43806 5012 43812 5024
rect 43767 4984 43812 5012
rect 43806 4972 43812 4984
rect 43864 4972 43870 5024
rect 44450 5012 44456 5024
rect 44411 4984 44456 5012
rect 44450 4972 44456 4984
rect 44508 4972 44514 5024
rect 46014 4972 46020 5024
rect 46072 5012 46078 5024
rect 47673 5015 47731 5021
rect 47673 5012 47685 5015
rect 46072 4984 47685 5012
rect 46072 4972 46078 4984
rect 47673 4981 47685 4984
rect 47719 4981 47731 5015
rect 47673 4975 47731 4981
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 3237 4811 3295 4817
rect 3237 4777 3249 4811
rect 3283 4808 3295 4811
rect 4062 4808 4068 4820
rect 3283 4780 4068 4808
rect 3283 4777 3295 4780
rect 3237 4771 3295 4777
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 31662 4768 31668 4820
rect 31720 4808 31726 4820
rect 32125 4811 32183 4817
rect 32125 4808 32137 4811
rect 31720 4780 32137 4808
rect 31720 4768 31726 4780
rect 32125 4777 32137 4780
rect 32171 4777 32183 4811
rect 32125 4771 32183 4777
rect 33229 4811 33287 4817
rect 33229 4777 33241 4811
rect 33275 4808 33287 4811
rect 33410 4808 33416 4820
rect 33275 4780 33416 4808
rect 33275 4777 33287 4780
rect 33229 4771 33287 4777
rect 33410 4768 33416 4780
rect 33468 4768 33474 4820
rect 44361 4811 44419 4817
rect 44361 4777 44373 4811
rect 44407 4808 44419 4811
rect 45646 4808 45652 4820
rect 44407 4780 45652 4808
rect 44407 4777 44419 4780
rect 44361 4771 44419 4777
rect 45646 4768 45652 4780
rect 45704 4768 45710 4820
rect 4890 4740 4896 4752
rect 3068 4712 4896 4740
rect 1673 4675 1731 4681
rect 1673 4641 1685 4675
rect 1719 4672 1731 4675
rect 2866 4672 2872 4684
rect 1719 4644 2872 4672
rect 1719 4641 1731 4644
rect 1673 4635 1731 4641
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4573 1639 4607
rect 1581 4567 1639 4573
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4573 1823 4607
rect 1765 4567 1823 4573
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4604 2283 4607
rect 2682 4604 2688 4616
rect 2271 4576 2688 4604
rect 2271 4573 2283 4576
rect 2225 4567 2283 4573
rect 1596 4468 1624 4567
rect 1780 4536 1808 4567
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 3068 4613 3096 4712
rect 4890 4700 4896 4712
rect 4948 4700 4954 4752
rect 10318 4740 10324 4752
rect 8956 4712 10324 4740
rect 3234 4632 3240 4684
rect 3292 4672 3298 4684
rect 3789 4675 3847 4681
rect 3789 4672 3801 4675
rect 3292 4644 3801 4672
rect 3292 4632 3298 4644
rect 3789 4641 3801 4644
rect 3835 4641 3847 4675
rect 4246 4672 4252 4684
rect 4207 4644 4252 4672
rect 3789 4635 3847 4641
rect 4246 4632 4252 4644
rect 4304 4632 4310 4684
rect 5534 4632 5540 4684
rect 5592 4672 5598 4684
rect 6178 4672 6184 4684
rect 5592 4644 6184 4672
rect 5592 4632 5598 4644
rect 6178 4632 6184 4644
rect 6236 4672 6242 4684
rect 6273 4675 6331 4681
rect 6273 4672 6285 4675
rect 6236 4644 6285 4672
rect 6236 4632 6242 4644
rect 6273 4641 6285 4644
rect 6319 4641 6331 4675
rect 6454 4672 6460 4684
rect 6415 4644 6460 4672
rect 6273 4635 6331 4641
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 6914 4672 6920 4684
rect 6875 4644 6920 4672
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 8956 4681 8984 4712
rect 10318 4700 10324 4712
rect 10376 4700 10382 4752
rect 14737 4743 14795 4749
rect 14737 4709 14749 4743
rect 14783 4740 14795 4743
rect 14918 4740 14924 4752
rect 14783 4712 14924 4740
rect 14783 4709 14795 4712
rect 14737 4703 14795 4709
rect 14918 4700 14924 4712
rect 14976 4700 14982 4752
rect 19797 4743 19855 4749
rect 19797 4709 19809 4743
rect 19843 4740 19855 4743
rect 24946 4740 24952 4752
rect 19843 4712 24952 4740
rect 19843 4709 19855 4712
rect 19797 4703 19855 4709
rect 24946 4700 24952 4712
rect 25004 4700 25010 4752
rect 34790 4740 34796 4752
rect 26206 4712 34796 4740
rect 8941 4675 8999 4681
rect 8941 4641 8953 4675
rect 8987 4641 8999 4675
rect 8941 4635 8999 4641
rect 9125 4675 9183 4681
rect 9125 4641 9137 4675
rect 9171 4672 9183 4675
rect 9214 4672 9220 4684
rect 9171 4644 9220 4672
rect 9171 4641 9183 4644
rect 9125 4635 9183 4641
rect 9214 4632 9220 4644
rect 9272 4632 9278 4684
rect 9766 4672 9772 4684
rect 9727 4644 9772 4672
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4672 11483 4675
rect 26206 4672 26234 4712
rect 34790 4700 34796 4712
rect 34848 4700 34854 4752
rect 11471 4644 26234 4672
rect 27341 4675 27399 4681
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 27341 4641 27353 4675
rect 27387 4672 27399 4675
rect 28902 4672 28908 4684
rect 27387 4644 28908 4672
rect 27387 4641 27399 4644
rect 27341 4635 27399 4641
rect 28902 4632 28908 4644
rect 28960 4632 28966 4684
rect 45830 4672 45836 4684
rect 35452 4644 36676 4672
rect 35452 4616 35480 4644
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4573 3111 4607
rect 3053 4567 3111 4573
rect 15289 4607 15347 4613
rect 15289 4573 15301 4607
rect 15335 4604 15347 4607
rect 15838 4604 15844 4616
rect 15335 4576 15844 4604
rect 15335 4573 15347 4576
rect 15289 4567 15347 4573
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 16114 4604 16120 4616
rect 16075 4576 16120 4604
rect 16114 4564 16120 4576
rect 16172 4564 16178 4616
rect 16758 4604 16764 4616
rect 16719 4576 16764 4604
rect 16758 4564 16764 4576
rect 16816 4564 16822 4616
rect 17126 4564 17132 4616
rect 17184 4604 17190 4616
rect 17405 4607 17463 4613
rect 17405 4604 17417 4607
rect 17184 4576 17417 4604
rect 17184 4564 17190 4576
rect 17405 4573 17417 4576
rect 17451 4573 17463 4607
rect 18046 4604 18052 4616
rect 18007 4576 18052 4604
rect 17405 4567 17463 4573
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 18414 4564 18420 4616
rect 18472 4604 18478 4616
rect 18509 4607 18567 4613
rect 18509 4604 18521 4607
rect 18472 4576 18521 4604
rect 18472 4564 18478 4576
rect 18509 4573 18521 4576
rect 18555 4573 18567 4607
rect 18509 4567 18567 4573
rect 20257 4607 20315 4613
rect 20257 4573 20269 4607
rect 20303 4573 20315 4607
rect 20530 4604 20536 4616
rect 20491 4576 20536 4604
rect 20257 4567 20315 4573
rect 2866 4536 2872 4548
rect 1780 4508 2872 4536
rect 2866 4496 2872 4508
rect 2924 4496 2930 4548
rect 3602 4496 3608 4548
rect 3660 4536 3666 4548
rect 3973 4539 4031 4545
rect 3973 4536 3985 4539
rect 3660 4508 3985 4536
rect 3660 4496 3666 4508
rect 3973 4505 3985 4508
rect 4019 4505 4031 4539
rect 3973 4499 4031 4505
rect 11609 4539 11667 4545
rect 11609 4505 11621 4539
rect 11655 4536 11667 4539
rect 12434 4536 12440 4548
rect 11655 4508 12440 4536
rect 11655 4505 11667 4508
rect 11609 4499 11667 4505
rect 12434 4496 12440 4508
rect 12492 4496 12498 4548
rect 13265 4539 13323 4545
rect 13265 4505 13277 4539
rect 13311 4536 13323 4539
rect 13630 4536 13636 4548
rect 13311 4508 13636 4536
rect 13311 4505 13323 4508
rect 13265 4499 13323 4505
rect 13630 4496 13636 4508
rect 13688 4496 13694 4548
rect 14553 4539 14611 4545
rect 14553 4505 14565 4539
rect 14599 4536 14611 4539
rect 14642 4536 14648 4548
rect 14599 4508 14648 4536
rect 14599 4505 14611 4508
rect 14553 4499 14611 4505
rect 14642 4496 14648 4508
rect 14700 4496 14706 4548
rect 19426 4496 19432 4548
rect 19484 4536 19490 4548
rect 19613 4539 19671 4545
rect 19613 4536 19625 4539
rect 19484 4508 19625 4536
rect 19484 4496 19490 4508
rect 19613 4505 19625 4508
rect 19659 4536 19671 4539
rect 20272 4536 20300 4567
rect 20530 4564 20536 4576
rect 20588 4564 20594 4616
rect 21910 4604 21916 4616
rect 21871 4576 21916 4604
rect 21910 4564 21916 4576
rect 21968 4564 21974 4616
rect 22373 4607 22431 4613
rect 22373 4573 22385 4607
rect 22419 4573 22431 4607
rect 22373 4567 22431 4573
rect 23017 4607 23075 4613
rect 23017 4573 23029 4607
rect 23063 4604 23075 4607
rect 23290 4604 23296 4616
rect 23063 4576 23296 4604
rect 23063 4573 23075 4576
rect 23017 4567 23075 4573
rect 19659 4508 20300 4536
rect 19659 4505 19671 4508
rect 19613 4499 19671 4505
rect 21082 4496 21088 4548
rect 21140 4536 21146 4548
rect 22388 4536 22416 4567
rect 23290 4564 23296 4576
rect 23348 4604 23354 4616
rect 23661 4607 23719 4613
rect 23661 4604 23673 4607
rect 23348 4576 23673 4604
rect 23348 4564 23354 4576
rect 23661 4573 23673 4576
rect 23707 4604 23719 4607
rect 24581 4607 24639 4613
rect 24581 4604 24593 4607
rect 23707 4576 24593 4604
rect 23707 4573 23719 4576
rect 23661 4567 23719 4573
rect 24581 4573 24593 4576
rect 24627 4604 24639 4607
rect 25225 4607 25283 4613
rect 25225 4604 25237 4607
rect 24627 4576 25237 4604
rect 24627 4573 24639 4576
rect 24581 4567 24639 4573
rect 25225 4573 25237 4576
rect 25271 4573 25283 4607
rect 25225 4567 25283 4573
rect 25314 4564 25320 4616
rect 25372 4604 25378 4616
rect 26053 4607 26111 4613
rect 26053 4604 26065 4607
rect 25372 4576 26065 4604
rect 25372 4564 25378 4576
rect 26053 4573 26065 4576
rect 26099 4573 26111 4607
rect 26053 4567 26111 4573
rect 27614 4564 27620 4616
rect 27672 4604 27678 4616
rect 28077 4607 28135 4613
rect 28077 4604 28089 4607
rect 27672 4576 28089 4604
rect 27672 4564 27678 4576
rect 28077 4573 28089 4576
rect 28123 4604 28135 4607
rect 28534 4604 28540 4616
rect 28123 4576 28540 4604
rect 28123 4573 28135 4576
rect 28077 4567 28135 4573
rect 28534 4564 28540 4576
rect 28592 4564 28598 4616
rect 29730 4604 29736 4616
rect 29691 4576 29736 4604
rect 29730 4564 29736 4576
rect 29788 4564 29794 4616
rect 30374 4604 30380 4616
rect 30335 4576 30380 4604
rect 30374 4564 30380 4576
rect 30432 4564 30438 4616
rect 31021 4607 31079 4613
rect 31021 4573 31033 4607
rect 31067 4604 31079 4607
rect 31754 4604 31760 4616
rect 31067 4576 31760 4604
rect 31067 4573 31079 4576
rect 31021 4567 31079 4573
rect 31754 4564 31760 4576
rect 31812 4564 31818 4616
rect 33965 4607 34023 4613
rect 33965 4573 33977 4607
rect 34011 4604 34023 4607
rect 34422 4604 34428 4616
rect 34011 4576 34428 4604
rect 34011 4573 34023 4576
rect 33965 4567 34023 4573
rect 34422 4564 34428 4576
rect 34480 4564 34486 4616
rect 34790 4564 34796 4616
rect 34848 4604 34854 4616
rect 34885 4607 34943 4613
rect 34885 4604 34897 4607
rect 34848 4576 34897 4604
rect 34848 4564 34854 4576
rect 34885 4573 34897 4576
rect 34931 4573 34943 4607
rect 34885 4567 34943 4573
rect 35345 4607 35403 4613
rect 35345 4573 35357 4607
rect 35391 4604 35403 4607
rect 35434 4604 35440 4616
rect 35391 4576 35440 4604
rect 35391 4573 35403 4576
rect 35345 4567 35403 4573
rect 35434 4564 35440 4576
rect 35492 4564 35498 4616
rect 36170 4604 36176 4616
rect 36131 4576 36176 4604
rect 36170 4564 36176 4576
rect 36228 4564 36234 4616
rect 36648 4613 36676 4644
rect 37568 4644 44312 4672
rect 45791 4644 45836 4672
rect 36633 4607 36691 4613
rect 36633 4573 36645 4607
rect 36679 4573 36691 4607
rect 36633 4567 36691 4573
rect 21140 4508 22416 4536
rect 21140 4496 21146 4508
rect 23382 4496 23388 4548
rect 23440 4536 23446 4548
rect 37568 4545 37596 4644
rect 37737 4607 37795 4613
rect 37737 4573 37749 4607
rect 37783 4604 37795 4607
rect 37918 4604 37924 4616
rect 37783 4576 37924 4604
rect 37783 4573 37795 4576
rect 37737 4567 37795 4573
rect 37918 4564 37924 4576
rect 37976 4604 37982 4616
rect 38197 4607 38255 4613
rect 38197 4604 38209 4607
rect 37976 4576 38209 4604
rect 37976 4564 37982 4576
rect 38197 4573 38209 4576
rect 38243 4573 38255 4607
rect 39022 4604 39028 4616
rect 38983 4576 39028 4604
rect 38197 4567 38255 4573
rect 27893 4539 27951 4545
rect 27893 4536 27905 4539
rect 23440 4508 27905 4536
rect 23440 4496 23446 4508
rect 27893 4505 27905 4508
rect 27939 4536 27951 4539
rect 32033 4539 32091 4545
rect 32033 4536 32045 4539
rect 27939 4508 32045 4536
rect 27939 4505 27951 4508
rect 27893 4499 27951 4505
rect 32033 4505 32045 4508
rect 32079 4536 32091 4539
rect 33137 4539 33195 4545
rect 33137 4536 33149 4539
rect 32079 4508 33149 4536
rect 32079 4505 32091 4508
rect 32033 4499 32091 4505
rect 33137 4505 33149 4508
rect 33183 4505 33195 4539
rect 33137 4499 33195 4505
rect 37553 4539 37611 4545
rect 37553 4505 37565 4539
rect 37599 4505 37611 4539
rect 38212 4536 38240 4567
rect 39022 4564 39028 4576
rect 39080 4564 39086 4616
rect 40788 4613 40816 4644
rect 39853 4607 39911 4613
rect 39853 4573 39865 4607
rect 39899 4573 39911 4607
rect 39853 4567 39911 4573
rect 40773 4607 40831 4613
rect 40773 4573 40785 4607
rect 40819 4573 40831 4607
rect 40773 4567 40831 4573
rect 40957 4607 41015 4613
rect 40957 4573 40969 4607
rect 41003 4604 41015 4607
rect 41417 4607 41475 4613
rect 41417 4604 41429 4607
rect 41003 4576 41429 4604
rect 41003 4573 41015 4576
rect 40957 4567 41015 4573
rect 41417 4573 41429 4576
rect 41463 4573 41475 4607
rect 42242 4604 42248 4616
rect 42203 4576 42248 4604
rect 41417 4567 41475 4573
rect 39868 4536 39896 4567
rect 38212 4508 39896 4536
rect 41432 4536 41460 4567
rect 42242 4564 42248 4576
rect 42300 4564 42306 4616
rect 42426 4564 42432 4616
rect 42484 4604 42490 4616
rect 42705 4607 42763 4613
rect 42705 4604 42717 4607
rect 42484 4576 42717 4604
rect 42484 4564 42490 4576
rect 42705 4573 42717 4576
rect 42751 4573 42763 4607
rect 43530 4604 43536 4616
rect 43491 4576 43536 4604
rect 42705 4567 42763 4573
rect 43530 4564 43536 4576
rect 43588 4564 43594 4616
rect 44284 4613 44312 4644
rect 45830 4632 45836 4644
rect 45888 4632 45894 4684
rect 46014 4672 46020 4684
rect 45975 4644 46020 4672
rect 46014 4632 46020 4644
rect 46072 4632 46078 4684
rect 46474 4672 46480 4684
rect 46435 4644 46480 4672
rect 46474 4632 46480 4644
rect 46532 4632 46538 4684
rect 44269 4607 44327 4613
rect 44269 4573 44281 4607
rect 44315 4604 44327 4607
rect 45189 4607 45247 4613
rect 45189 4604 45201 4607
rect 44315 4576 45201 4604
rect 44315 4573 44327 4576
rect 44269 4567 44327 4573
rect 45189 4573 45201 4576
rect 45235 4573 45247 4607
rect 45189 4567 45247 4573
rect 42444 4536 42472 4564
rect 41432 4508 42472 4536
rect 37553 4499 37611 4505
rect 2222 4468 2228 4480
rect 1596 4440 2228 4468
rect 2222 4428 2228 4440
rect 2280 4428 2286 4480
rect 2317 4471 2375 4477
rect 2317 4437 2329 4471
rect 2363 4468 2375 4471
rect 6454 4468 6460 4480
rect 2363 4440 6460 4468
rect 2363 4437 2375 4440
rect 2317 4431 2375 4437
rect 6454 4428 6460 4440
rect 6512 4428 6518 4480
rect 15378 4468 15384 4480
rect 15339 4440 15384 4468
rect 15378 4428 15384 4440
rect 15436 4428 15442 4480
rect 18601 4471 18659 4477
rect 18601 4437 18613 4471
rect 18647 4468 18659 4471
rect 18690 4468 18696 4480
rect 18647 4440 18696 4468
rect 18647 4437 18659 4440
rect 18601 4431 18659 4437
rect 18690 4428 18696 4440
rect 18748 4428 18754 4480
rect 22094 4428 22100 4480
rect 22152 4468 22158 4480
rect 22465 4471 22523 4477
rect 22465 4468 22477 4471
rect 22152 4440 22477 4468
rect 22152 4428 22158 4440
rect 22465 4437 22477 4440
rect 22511 4437 22523 4471
rect 23106 4468 23112 4480
rect 23067 4440 23112 4468
rect 22465 4431 22523 4437
rect 23106 4428 23112 4440
rect 23164 4428 23170 4480
rect 23753 4471 23811 4477
rect 23753 4437 23765 4471
rect 23799 4468 23811 4471
rect 24026 4468 24032 4480
rect 23799 4440 24032 4468
rect 23799 4437 23811 4440
rect 23753 4431 23811 4437
rect 24026 4428 24032 4440
rect 24084 4428 24090 4480
rect 24673 4471 24731 4477
rect 24673 4437 24685 4471
rect 24719 4468 24731 4471
rect 24762 4468 24768 4480
rect 24719 4440 24768 4468
rect 24719 4437 24731 4440
rect 24673 4431 24731 4437
rect 24762 4428 24768 4440
rect 24820 4428 24826 4480
rect 25317 4471 25375 4477
rect 25317 4437 25329 4471
rect 25363 4468 25375 4471
rect 25866 4468 25872 4480
rect 25363 4440 25872 4468
rect 25363 4437 25375 4440
rect 25317 4431 25375 4437
rect 25866 4428 25872 4440
rect 25924 4428 25930 4480
rect 28629 4471 28687 4477
rect 28629 4437 28641 4471
rect 28675 4468 28687 4471
rect 29454 4468 29460 4480
rect 28675 4440 29460 4468
rect 28675 4437 28687 4440
rect 28629 4431 28687 4437
rect 29454 4428 29460 4440
rect 29512 4428 29518 4480
rect 35434 4468 35440 4480
rect 35395 4440 35440 4468
rect 35434 4428 35440 4440
rect 35492 4428 35498 4480
rect 36725 4471 36783 4477
rect 36725 4437 36737 4471
rect 36771 4468 36783 4471
rect 37458 4468 37464 4480
rect 36771 4440 37464 4468
rect 36771 4437 36783 4440
rect 36725 4431 36783 4437
rect 37458 4428 37464 4440
rect 37516 4428 37522 4480
rect 37568 4468 37596 4499
rect 45002 4496 45008 4548
rect 45060 4536 45066 4548
rect 45370 4536 45376 4548
rect 45060 4508 45376 4536
rect 45060 4496 45066 4508
rect 45370 4496 45376 4508
rect 45428 4496 45434 4548
rect 37734 4468 37740 4480
rect 37568 4440 37740 4468
rect 37734 4428 37740 4440
rect 37792 4428 37798 4480
rect 38286 4468 38292 4480
rect 38247 4440 38292 4468
rect 38286 4428 38292 4440
rect 38344 4428 38350 4480
rect 39945 4471 40003 4477
rect 39945 4437 39957 4471
rect 39991 4468 40003 4471
rect 40034 4468 40040 4480
rect 39991 4440 40040 4468
rect 39991 4437 40003 4440
rect 39945 4431 40003 4437
rect 40034 4428 40040 4440
rect 40092 4428 40098 4480
rect 41506 4468 41512 4480
rect 41467 4440 41512 4468
rect 41506 4428 41512 4440
rect 41564 4428 41570 4480
rect 42794 4468 42800 4480
rect 42755 4440 42800 4468
rect 42794 4428 42800 4440
rect 42852 4428 42858 4480
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 2222 4224 2228 4276
rect 2280 4264 2286 4276
rect 5534 4264 5540 4276
rect 2280 4236 5540 4264
rect 2280 4224 2286 4236
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 20530 4224 20536 4276
rect 20588 4264 20594 4276
rect 23290 4264 23296 4276
rect 20588 4236 23152 4264
rect 23251 4236 23296 4264
rect 20588 4224 20594 4236
rect 2314 4156 2320 4208
rect 2372 4196 2378 4208
rect 13906 4196 13912 4208
rect 2372 4168 12480 4196
rect 2372 4156 2378 4168
rect 1578 4128 1584 4140
rect 1539 4100 1584 4128
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 3970 4128 3976 4140
rect 3931 4100 3976 4128
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 1762 4060 1768 4072
rect 1723 4032 1768 4060
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 2041 4063 2099 4069
rect 2041 4029 2053 4063
rect 2087 4029 2099 4063
rect 2041 4023 2099 4029
rect 750 3952 756 4004
rect 808 3992 814 4004
rect 2056 3992 2084 4023
rect 3786 4020 3792 4072
rect 3844 4060 3850 4072
rect 4157 4063 4215 4069
rect 4157 4060 4169 4063
rect 3844 4032 4169 4060
rect 3844 4020 3850 4032
rect 4157 4029 4169 4032
rect 4203 4029 4215 4063
rect 4157 4023 4215 4029
rect 4433 4063 4491 4069
rect 4433 4029 4445 4063
rect 4479 4029 4491 4063
rect 4433 4023 4491 4029
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4029 6883 4063
rect 7006 4060 7012 4072
rect 6967 4032 7012 4060
rect 6825 4023 6883 4029
rect 808 3964 2084 3992
rect 808 3952 814 3964
rect 3326 3952 3332 4004
rect 3384 3992 3390 4004
rect 4246 3992 4252 4004
rect 3384 3964 4252 3992
rect 3384 3952 3390 3964
rect 4246 3952 4252 3964
rect 4304 3952 4310 4004
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 4448 3924 4476 4023
rect 6840 3992 6868 4023
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 7190 4020 7196 4072
rect 7248 4060 7254 4072
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 7248 4032 7297 4060
rect 7248 4020 7254 4032
rect 7285 4029 7297 4032
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4029 9183 4063
rect 9306 4060 9312 4072
rect 9267 4032 9312 4060
rect 9125 4023 9183 4029
rect 7098 3992 7104 4004
rect 6840 3964 7104 3992
rect 7098 3952 7104 3964
rect 7156 3952 7162 4004
rect 9140 3992 9168 4023
rect 9306 4020 9312 4032
rect 9364 4020 9370 4072
rect 10965 4063 11023 4069
rect 10965 4029 10977 4063
rect 11011 4060 11023 4063
rect 11698 4060 11704 4072
rect 11011 4032 11704 4060
rect 11011 4029 11023 4032
rect 10965 4023 11023 4029
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 12452 4060 12480 4168
rect 13280 4168 13912 4196
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4128 12587 4131
rect 13280 4128 13308 4168
rect 13906 4156 13912 4168
rect 13964 4196 13970 4208
rect 14642 4196 14648 4208
rect 13964 4168 14648 4196
rect 13964 4156 13970 4168
rect 14642 4156 14648 4168
rect 14700 4196 14706 4208
rect 15657 4199 15715 4205
rect 15657 4196 15669 4199
rect 14700 4168 15669 4196
rect 14700 4156 14706 4168
rect 15657 4165 15669 4168
rect 15703 4165 15715 4199
rect 18414 4196 18420 4208
rect 15657 4159 15715 4165
rect 17972 4168 18420 4196
rect 12575 4100 13308 4128
rect 12575 4097 12587 4100
rect 12529 4091 12587 4097
rect 15838 4088 15844 4140
rect 15896 4128 15902 4140
rect 16482 4128 16488 4140
rect 15896 4100 16488 4128
rect 15896 4088 15902 4100
rect 16482 4088 16488 4100
rect 16540 4128 16546 4140
rect 17221 4131 17279 4137
rect 17221 4128 17233 4131
rect 16540 4100 17233 4128
rect 16540 4088 16546 4100
rect 17221 4097 17233 4100
rect 17267 4097 17279 4131
rect 17221 4091 17279 4097
rect 17865 4131 17923 4137
rect 17865 4097 17877 4131
rect 17911 4128 17923 4131
rect 17972 4128 18000 4168
rect 18414 4156 18420 4168
rect 18472 4156 18478 4208
rect 18690 4196 18696 4208
rect 18651 4168 18696 4196
rect 18690 4156 18696 4168
rect 18748 4156 18754 4208
rect 20916 4205 20944 4236
rect 20901 4199 20959 4205
rect 20901 4165 20913 4199
rect 20947 4165 20959 4199
rect 21082 4196 21088 4208
rect 21043 4168 21088 4196
rect 20901 4159 20959 4165
rect 21082 4156 21088 4168
rect 21140 4156 21146 4208
rect 17911 4100 18000 4128
rect 17911 4097 17923 4100
rect 17865 4091 17923 4097
rect 18046 4088 18052 4140
rect 18104 4128 18110 4140
rect 18509 4131 18567 4137
rect 18509 4128 18521 4131
rect 18104 4100 18521 4128
rect 18104 4088 18110 4100
rect 18509 4097 18521 4100
rect 18555 4097 18567 4131
rect 18509 4091 18567 4097
rect 22465 4131 22523 4137
rect 22465 4097 22477 4131
rect 22511 4097 22523 4131
rect 23124 4128 23152 4236
rect 23290 4224 23296 4236
rect 23348 4224 23354 4276
rect 23382 4156 23388 4208
rect 23440 4156 23446 4208
rect 24026 4196 24032 4208
rect 23987 4168 24032 4196
rect 24026 4156 24032 4168
rect 24084 4156 24090 4208
rect 28442 4196 28448 4208
rect 28403 4168 28448 4196
rect 28442 4156 28448 4168
rect 28500 4156 28506 4208
rect 32306 4196 32312 4208
rect 32267 4168 32312 4196
rect 32306 4156 32312 4168
rect 32364 4156 32370 4208
rect 34885 4199 34943 4205
rect 34885 4165 34897 4199
rect 34931 4196 34943 4199
rect 35342 4196 35348 4208
rect 34931 4168 35348 4196
rect 34931 4165 34943 4168
rect 34885 4159 34943 4165
rect 35342 4156 35348 4168
rect 35400 4156 35406 4208
rect 37550 4196 37556 4208
rect 37511 4168 37556 4196
rect 37550 4156 37556 4168
rect 37608 4156 37614 4208
rect 43254 4196 43260 4208
rect 42628 4168 43260 4196
rect 23201 4131 23259 4137
rect 23201 4128 23213 4131
rect 23124 4100 23213 4128
rect 22465 4091 22523 4097
rect 23201 4097 23213 4100
rect 23247 4128 23259 4131
rect 23400 4128 23428 4156
rect 23842 4128 23848 4140
rect 23247 4100 23428 4128
rect 23803 4100 23848 4128
rect 23247 4097 23259 4100
rect 23201 4091 23259 4097
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12452 4032 12817 4060
rect 12805 4029 12817 4032
rect 12851 4060 12863 4063
rect 13078 4060 13084 4072
rect 12851 4032 13084 4060
rect 12851 4029 12863 4032
rect 12805 4023 12863 4029
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 13262 4060 13268 4072
rect 13223 4032 13268 4060
rect 13262 4020 13268 4032
rect 13320 4020 13326 4072
rect 13446 4060 13452 4072
rect 13407 4032 13452 4060
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 15105 4063 15163 4069
rect 15105 4029 15117 4063
rect 15151 4060 15163 4063
rect 15562 4060 15568 4072
rect 15151 4032 15568 4060
rect 15151 4029 15163 4032
rect 15105 4023 15163 4029
rect 15562 4020 15568 4032
rect 15620 4020 15626 4072
rect 20070 4060 20076 4072
rect 20031 4032 20076 4060
rect 20070 4020 20076 4032
rect 20128 4020 20134 4072
rect 22480 4060 22508 4091
rect 23842 4088 23848 4100
rect 23900 4088 23906 4140
rect 27614 4128 27620 4140
rect 27575 4100 27620 4128
rect 27614 4088 27620 4100
rect 27672 4088 27678 4140
rect 31205 4131 31263 4137
rect 31205 4097 31217 4131
rect 31251 4128 31263 4131
rect 31662 4128 31668 4140
rect 31251 4100 31668 4128
rect 31251 4097 31263 4100
rect 31205 4091 31263 4097
rect 31662 4088 31668 4100
rect 31720 4088 31726 4140
rect 32122 4128 32128 4140
rect 32083 4100 32128 4128
rect 32122 4088 32128 4100
rect 32180 4088 32186 4140
rect 42628 4137 42656 4168
rect 43254 4156 43260 4168
rect 43312 4156 43318 4208
rect 42613 4131 42671 4137
rect 42613 4097 42625 4131
rect 42659 4097 42671 4131
rect 42613 4091 42671 4097
rect 23290 4060 23296 4072
rect 22480 4032 23296 4060
rect 23290 4020 23296 4032
rect 23348 4020 23354 4072
rect 24486 4060 24492 4072
rect 24447 4032 24492 4060
rect 24486 4020 24492 4032
rect 24544 4020 24550 4072
rect 28261 4063 28319 4069
rect 28261 4029 28273 4063
rect 28307 4060 28319 4063
rect 29730 4060 29736 4072
rect 28307 4032 29736 4060
rect 28307 4029 28319 4032
rect 28261 4023 28319 4029
rect 29730 4020 29736 4032
rect 29788 4020 29794 4072
rect 29825 4063 29883 4069
rect 29825 4029 29837 4063
rect 29871 4029 29883 4063
rect 32950 4060 32956 4072
rect 32911 4032 32956 4060
rect 29825 4023 29883 4029
rect 25222 3992 25228 4004
rect 9140 3964 25228 3992
rect 25222 3952 25228 3964
rect 25280 3952 25286 4004
rect 26234 3952 26240 4004
rect 26292 3992 26298 4004
rect 26292 3964 27844 3992
rect 26292 3952 26298 3964
rect 4028 3896 4476 3924
rect 4028 3884 4034 3896
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 16298 3924 16304 3936
rect 13136 3896 16304 3924
rect 13136 3884 13142 3896
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 17034 3884 17040 3936
rect 17092 3924 17098 3936
rect 17313 3927 17371 3933
rect 17313 3924 17325 3927
rect 17092 3896 17325 3924
rect 17092 3884 17098 3896
rect 17313 3893 17325 3896
rect 17359 3893 17371 3927
rect 17313 3887 17371 3893
rect 17957 3927 18015 3933
rect 17957 3893 17969 3927
rect 18003 3924 18015 3927
rect 19426 3924 19432 3936
rect 18003 3896 19432 3924
rect 18003 3893 18015 3896
rect 17957 3887 18015 3893
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 22002 3924 22008 3936
rect 21963 3896 22008 3924
rect 22002 3884 22008 3896
rect 22060 3884 22066 3936
rect 22462 3884 22468 3936
rect 22520 3924 22526 3936
rect 22557 3927 22615 3933
rect 22557 3924 22569 3927
rect 22520 3896 22569 3924
rect 22520 3884 22526 3896
rect 22557 3893 22569 3896
rect 22603 3893 22615 3927
rect 22557 3887 22615 3893
rect 25682 3884 25688 3936
rect 25740 3924 25746 3936
rect 26329 3927 26387 3933
rect 26329 3924 26341 3927
rect 25740 3896 26341 3924
rect 25740 3884 25746 3896
rect 26329 3893 26341 3896
rect 26375 3893 26387 3927
rect 26329 3887 26387 3893
rect 26970 3884 26976 3936
rect 27028 3924 27034 3936
rect 27157 3927 27215 3933
rect 27157 3924 27169 3927
rect 27028 3896 27169 3924
rect 27028 3884 27034 3896
rect 27157 3893 27169 3896
rect 27203 3893 27215 3927
rect 27157 3887 27215 3893
rect 27614 3884 27620 3936
rect 27672 3924 27678 3936
rect 27709 3927 27767 3933
rect 27709 3924 27721 3927
rect 27672 3896 27721 3924
rect 27672 3884 27678 3896
rect 27709 3893 27721 3896
rect 27755 3893 27767 3927
rect 27816 3924 27844 3964
rect 29178 3952 29184 4004
rect 29236 3992 29242 4004
rect 29840 3992 29868 4023
rect 32950 4020 32956 4032
rect 33008 4020 33014 4072
rect 34701 4063 34759 4069
rect 34701 4029 34713 4063
rect 34747 4029 34759 4063
rect 36170 4060 36176 4072
rect 34701 4023 34759 4029
rect 35268 4032 36176 4060
rect 32490 3992 32496 4004
rect 29236 3964 29868 3992
rect 29932 3964 32496 3992
rect 29236 3952 29242 3964
rect 29932 3924 29960 3964
rect 32490 3952 32496 3964
rect 32548 3952 32554 4004
rect 34716 3992 34744 4023
rect 35268 3992 35296 4032
rect 36170 4020 36176 4032
rect 36228 4020 36234 4072
rect 36265 4063 36323 4069
rect 36265 4029 36277 4063
rect 36311 4029 36323 4063
rect 36265 4023 36323 4029
rect 37369 4063 37427 4069
rect 37369 4029 37381 4063
rect 37415 4029 37427 4063
rect 38102 4060 38108 4072
rect 38063 4032 38108 4060
rect 37369 4023 37427 4029
rect 34716 3964 35296 3992
rect 35526 3952 35532 4004
rect 35584 3992 35590 4004
rect 36280 3992 36308 4023
rect 35584 3964 36308 3992
rect 37384 3992 37412 4023
rect 38102 4020 38108 4032
rect 38160 4020 38166 4072
rect 40037 4063 40095 4069
rect 40037 4029 40049 4063
rect 40083 4029 40095 4063
rect 40037 4023 40095 4029
rect 40221 4063 40279 4069
rect 40221 4029 40233 4063
rect 40267 4060 40279 4063
rect 41506 4060 41512 4072
rect 40267 4032 41512 4060
rect 40267 4029 40279 4032
rect 40221 4023 40279 4029
rect 39022 3992 39028 4004
rect 37384 3964 39028 3992
rect 35584 3952 35590 3964
rect 39022 3952 39028 3964
rect 39080 3952 39086 4004
rect 40052 3992 40080 4023
rect 41506 4020 41512 4032
rect 41564 4020 41570 4072
rect 41601 4063 41659 4069
rect 41601 4029 41613 4063
rect 41647 4029 41659 4063
rect 41601 4023 41659 4029
rect 42797 4063 42855 4069
rect 42797 4029 42809 4063
rect 42843 4060 42855 4063
rect 43806 4060 43812 4072
rect 42843 4032 43812 4060
rect 42843 4029 42855 4032
rect 42797 4023 42855 4029
rect 40126 3992 40132 4004
rect 40052 3964 40132 3992
rect 40126 3952 40132 3964
rect 40184 3952 40190 4004
rect 40678 3952 40684 4004
rect 40736 3992 40742 4004
rect 41616 3992 41644 4023
rect 43806 4020 43812 4032
rect 43864 4020 43870 4072
rect 43993 4063 44051 4069
rect 43993 4029 44005 4063
rect 44039 4029 44051 4063
rect 43993 4023 44051 4029
rect 45005 4063 45063 4069
rect 45005 4029 45017 4063
rect 45051 4029 45063 4063
rect 45186 4060 45192 4072
rect 45147 4032 45192 4060
rect 45005 4023 45063 4029
rect 40736 3964 41644 3992
rect 40736 3952 40742 3964
rect 43254 3952 43260 4004
rect 43312 3992 43318 4004
rect 44008 3992 44036 4023
rect 43312 3964 44036 3992
rect 45020 3992 45048 4023
rect 45186 4020 45192 4032
rect 45244 4020 45250 4072
rect 45830 4060 45836 4072
rect 45791 4032 45836 4060
rect 45830 4020 45836 4032
rect 45888 4020 45894 4072
rect 47765 3995 47823 4001
rect 47765 3992 47777 3995
rect 45020 3964 47777 3992
rect 43312 3952 43318 3964
rect 47765 3961 47777 3964
rect 47811 3961 47823 3995
rect 47765 3955 47823 3961
rect 30742 3924 30748 3936
rect 27816 3896 29960 3924
rect 30703 3896 30748 3924
rect 27709 3887 27767 3893
rect 30742 3884 30748 3896
rect 30800 3884 30806 3936
rect 31294 3924 31300 3936
rect 31255 3896 31300 3924
rect 31294 3884 31300 3896
rect 31352 3884 31358 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 1854 3720 1860 3732
rect 1412 3692 1860 3720
rect 1412 3593 1440 3692
rect 1854 3680 1860 3692
rect 1912 3680 1918 3732
rect 13262 3680 13268 3732
rect 13320 3720 13326 3732
rect 13320 3692 43484 3720
rect 13320 3680 13326 3692
rect 2866 3612 2872 3664
rect 2924 3652 2930 3664
rect 4982 3652 4988 3664
rect 2924 3624 4988 3652
rect 2924 3612 2930 3624
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 1578 3544 1584 3596
rect 1636 3584 1642 3596
rect 4264 3593 4292 3624
rect 4982 3612 4988 3624
rect 5040 3612 5046 3664
rect 9490 3652 9496 3664
rect 6564 3624 9496 3652
rect 1857 3587 1915 3593
rect 1857 3584 1869 3587
rect 1636 3556 1869 3584
rect 1636 3544 1642 3556
rect 1857 3553 1869 3556
rect 1903 3553 1915 3587
rect 1857 3547 1915 3553
rect 4249 3587 4307 3593
rect 4249 3553 4261 3587
rect 4295 3553 4307 3587
rect 4249 3547 4307 3553
rect 4433 3587 4491 3593
rect 4433 3553 4445 3587
rect 4479 3584 4491 3587
rect 5166 3584 5172 3596
rect 4479 3556 5172 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 5902 3584 5908 3596
rect 5863 3556 5908 3584
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 6564 3593 6592 3624
rect 9490 3612 9496 3624
rect 9548 3612 9554 3664
rect 12406 3624 22048 3652
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3553 6607 3587
rect 6549 3547 6607 3553
rect 8941 3587 8999 3593
rect 8941 3553 8953 3587
rect 8987 3584 8999 3587
rect 9582 3584 9588 3596
rect 8987 3556 9588 3584
rect 8987 3553 8999 3556
rect 8941 3547 8999 3553
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 10410 3584 10416 3596
rect 10371 3556 10416 3584
rect 10410 3544 10416 3556
rect 10468 3544 10474 3596
rect 11241 3587 11299 3593
rect 11241 3553 11253 3587
rect 11287 3584 11299 3587
rect 12406 3584 12434 3624
rect 11287 3556 12434 3584
rect 14185 3587 14243 3593
rect 11287 3553 11299 3556
rect 11241 3547 11299 3553
rect 14185 3553 14197 3587
rect 14231 3584 14243 3587
rect 14366 3584 14372 3596
rect 14231 3556 14372 3584
rect 14231 3553 14243 3556
rect 14185 3547 14243 3553
rect 14366 3544 14372 3556
rect 14424 3544 14430 3596
rect 16114 3544 16120 3596
rect 16172 3584 16178 3596
rect 16485 3587 16543 3593
rect 16485 3584 16497 3587
rect 16172 3556 16497 3584
rect 16172 3544 16178 3556
rect 16485 3553 16497 3556
rect 16531 3553 16543 3587
rect 16485 3547 16543 3553
rect 16669 3587 16727 3593
rect 16669 3553 16681 3587
rect 16715 3584 16727 3587
rect 17402 3584 17408 3596
rect 16715 3556 17408 3584
rect 16715 3553 16727 3556
rect 16669 3547 16727 3553
rect 17402 3544 17408 3556
rect 17460 3544 17466 3596
rect 18138 3584 18144 3596
rect 18099 3556 18144 3584
rect 18138 3544 18144 3556
rect 18196 3544 18202 3596
rect 19150 3544 19156 3596
rect 19208 3584 19214 3596
rect 19245 3587 19303 3593
rect 19245 3584 19257 3587
rect 19208 3556 19257 3584
rect 19208 3544 19214 3556
rect 19245 3553 19257 3556
rect 19291 3553 19303 3587
rect 19426 3584 19432 3596
rect 19387 3556 19432 3584
rect 19245 3547 19303 3553
rect 19426 3544 19432 3556
rect 19484 3544 19490 3596
rect 20714 3584 20720 3596
rect 20675 3556 20720 3584
rect 20714 3544 20720 3556
rect 20772 3544 20778 3596
rect 21637 3587 21695 3593
rect 21637 3553 21649 3587
rect 21683 3584 21695 3587
rect 21910 3584 21916 3596
rect 21683 3556 21916 3584
rect 21683 3553 21695 3556
rect 21637 3547 21695 3553
rect 21910 3544 21916 3556
rect 21968 3544 21974 3596
rect 22020 3584 22048 3624
rect 24946 3612 24952 3664
rect 25004 3652 25010 3664
rect 30374 3652 30380 3664
rect 25004 3624 29500 3652
rect 25004 3612 25010 3624
rect 26234 3584 26240 3596
rect 22020 3556 26240 3584
rect 26234 3544 26240 3556
rect 26292 3544 26298 3596
rect 26510 3584 26516 3596
rect 26471 3556 26516 3584
rect 26510 3544 26516 3556
rect 26568 3544 26574 3596
rect 24946 3516 24952 3528
rect 24907 3488 24952 3516
rect 24946 3476 24952 3488
rect 25004 3476 25010 3528
rect 25682 3516 25688 3528
rect 25643 3488 25688 3516
rect 25682 3476 25688 3488
rect 25740 3476 25746 3528
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 27985 3519 28043 3525
rect 27985 3516 27997 3519
rect 27764 3488 27997 3516
rect 27764 3476 27770 3488
rect 27985 3485 27997 3488
rect 28031 3485 28043 3519
rect 28810 3516 28816 3528
rect 28771 3488 28816 3516
rect 27985 3479 28043 3485
rect 28810 3476 28816 3488
rect 28868 3476 28874 3528
rect 1581 3451 1639 3457
rect 1581 3417 1593 3451
rect 1627 3448 1639 3451
rect 2038 3448 2044 3460
rect 1627 3420 2044 3448
rect 1627 3417 1639 3420
rect 1581 3411 1639 3417
rect 2038 3408 2044 3420
rect 2096 3408 2102 3460
rect 6270 3408 6276 3460
rect 6328 3448 6334 3460
rect 6733 3451 6791 3457
rect 6733 3448 6745 3451
rect 6328 3420 6745 3448
rect 6328 3408 6334 3420
rect 6733 3417 6745 3420
rect 6779 3417 6791 3451
rect 6733 3411 6791 3417
rect 8389 3451 8447 3457
rect 8389 3417 8401 3451
rect 8435 3448 8447 3451
rect 8478 3448 8484 3460
rect 8435 3420 8484 3448
rect 8435 3417 8447 3420
rect 8389 3411 8447 3417
rect 8478 3408 8484 3420
rect 8536 3408 8542 3460
rect 9125 3451 9183 3457
rect 9125 3417 9137 3451
rect 9171 3448 9183 3451
rect 11146 3448 11152 3460
rect 9171 3420 11152 3448
rect 9171 3417 9183 3420
rect 9125 3411 9183 3417
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 11422 3448 11428 3460
rect 11383 3420 11428 3448
rect 11422 3408 11428 3420
rect 11480 3408 11486 3460
rect 12986 3408 12992 3460
rect 13044 3448 13050 3460
rect 13081 3451 13139 3457
rect 13081 3448 13093 3451
rect 13044 3420 13093 3448
rect 13044 3408 13050 3420
rect 13081 3417 13093 3420
rect 13127 3417 13139 3451
rect 13081 3411 13139 3417
rect 14369 3451 14427 3457
rect 14369 3417 14381 3451
rect 14415 3448 14427 3451
rect 14458 3448 14464 3460
rect 14415 3420 14464 3448
rect 14415 3417 14427 3420
rect 14369 3411 14427 3417
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 16025 3451 16083 3457
rect 16025 3417 16037 3451
rect 16071 3448 16083 3451
rect 16206 3448 16212 3460
rect 16071 3420 16212 3448
rect 16071 3417 16083 3420
rect 16025 3411 16083 3417
rect 16206 3408 16212 3420
rect 16264 3408 16270 3460
rect 16298 3408 16304 3460
rect 16356 3448 16362 3460
rect 19518 3448 19524 3460
rect 16356 3420 19524 3448
rect 16356 3408 16362 3420
rect 19518 3408 19524 3420
rect 19576 3408 19582 3460
rect 21821 3451 21879 3457
rect 21821 3417 21833 3451
rect 21867 3448 21879 3451
rect 22094 3448 22100 3460
rect 21867 3420 22100 3448
rect 21867 3417 21879 3420
rect 21821 3411 21879 3417
rect 22094 3408 22100 3420
rect 22152 3408 22158 3460
rect 22646 3408 22652 3460
rect 22704 3448 22710 3460
rect 23477 3451 23535 3457
rect 23477 3448 23489 3451
rect 22704 3420 23489 3448
rect 22704 3408 22710 3420
rect 23477 3417 23489 3420
rect 23523 3417 23535 3451
rect 25866 3448 25872 3460
rect 25827 3420 25872 3448
rect 23477 3411 23535 3417
rect 25866 3408 25872 3420
rect 25924 3408 25930 3460
rect 14182 3340 14188 3392
rect 14240 3380 14246 3392
rect 15930 3380 15936 3392
rect 14240 3352 15936 3380
rect 14240 3340 14246 3352
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 16666 3340 16672 3392
rect 16724 3380 16730 3392
rect 21726 3380 21732 3392
rect 16724 3352 21732 3380
rect 16724 3340 16730 3352
rect 21726 3340 21732 3352
rect 21784 3340 21790 3392
rect 25038 3380 25044 3392
rect 24999 3352 25044 3380
rect 25038 3340 25044 3352
rect 25096 3340 25102 3392
rect 27154 3340 27160 3392
rect 27212 3380 27218 3392
rect 28077 3383 28135 3389
rect 28077 3380 28089 3383
rect 27212 3352 28089 3380
rect 27212 3340 27218 3352
rect 28077 3349 28089 3352
rect 28123 3349 28135 3383
rect 29472 3380 29500 3624
rect 29564 3624 30380 3652
rect 29564 3593 29592 3624
rect 30374 3612 30380 3624
rect 30432 3612 30438 3664
rect 31662 3612 31668 3664
rect 31720 3652 31726 3664
rect 31720 3624 32352 3652
rect 31720 3612 31726 3624
rect 29549 3587 29607 3593
rect 29549 3553 29561 3587
rect 29595 3553 29607 3587
rect 29549 3547 29607 3553
rect 29733 3587 29791 3593
rect 29733 3553 29745 3587
rect 29779 3584 29791 3587
rect 31294 3584 31300 3596
rect 29779 3556 31300 3584
rect 29779 3553 29791 3556
rect 29733 3547 29791 3553
rect 31294 3544 31300 3556
rect 31352 3544 31358 3596
rect 31846 3584 31852 3596
rect 31807 3556 31852 3584
rect 31846 3544 31852 3556
rect 31904 3544 31910 3596
rect 32030 3584 32036 3596
rect 31991 3556 32036 3584
rect 32030 3544 32036 3556
rect 32088 3544 32094 3596
rect 32324 3593 32352 3624
rect 36814 3612 36820 3664
rect 36872 3652 36878 3664
rect 36872 3624 37504 3652
rect 36872 3612 36878 3624
rect 32309 3587 32367 3593
rect 32309 3553 32321 3587
rect 32355 3553 32367 3587
rect 34698 3584 34704 3596
rect 34659 3556 34704 3584
rect 32309 3547 32367 3553
rect 34698 3544 34704 3556
rect 34756 3544 34762 3596
rect 34882 3544 34888 3596
rect 34940 3584 34946 3596
rect 35161 3587 35219 3593
rect 35161 3584 35173 3587
rect 34940 3556 35173 3584
rect 34940 3544 34946 3556
rect 35161 3553 35173 3556
rect 35207 3553 35219 3587
rect 35161 3547 35219 3553
rect 36354 3544 36360 3596
rect 36412 3584 36418 3596
rect 37001 3587 37059 3593
rect 37001 3584 37013 3587
rect 36412 3556 37013 3584
rect 36412 3544 36418 3556
rect 37001 3553 37013 3556
rect 37047 3553 37059 3587
rect 37001 3547 37059 3553
rect 37185 3587 37243 3593
rect 37185 3553 37197 3587
rect 37231 3584 37243 3587
rect 37366 3584 37372 3596
rect 37231 3556 37372 3584
rect 37231 3553 37243 3556
rect 37185 3547 37243 3553
rect 37366 3544 37372 3556
rect 37424 3544 37430 3596
rect 37476 3593 37504 3624
rect 40126 3612 40132 3664
rect 40184 3652 40190 3664
rect 40184 3624 40356 3652
rect 40184 3612 40190 3624
rect 37461 3587 37519 3593
rect 37461 3553 37473 3587
rect 37507 3553 37519 3587
rect 37461 3547 37519 3553
rect 39853 3587 39911 3593
rect 39853 3553 39865 3587
rect 39899 3584 39911 3587
rect 40218 3584 40224 3596
rect 39899 3556 40224 3584
rect 39899 3553 39911 3556
rect 39853 3547 39911 3553
rect 40218 3544 40224 3556
rect 40276 3544 40282 3596
rect 40328 3593 40356 3624
rect 41966 3612 41972 3664
rect 42024 3652 42030 3664
rect 43456 3652 43484 3692
rect 45370 3680 45376 3732
rect 45428 3720 45434 3732
rect 45428 3692 48176 3720
rect 45428 3680 45434 3692
rect 45554 3652 45560 3664
rect 42024 3624 42932 3652
rect 43456 3624 45560 3652
rect 42024 3612 42030 3624
rect 40313 3587 40371 3593
rect 40313 3553 40325 3587
rect 40359 3553 40371 3587
rect 40313 3547 40371 3553
rect 41598 3544 41604 3596
rect 41656 3584 41662 3596
rect 42153 3587 42211 3593
rect 42153 3584 42165 3587
rect 41656 3556 42165 3584
rect 41656 3544 41662 3556
rect 42153 3553 42165 3556
rect 42199 3553 42211 3587
rect 42153 3547 42211 3553
rect 42337 3587 42395 3593
rect 42337 3553 42349 3587
rect 42383 3584 42395 3587
rect 42794 3584 42800 3596
rect 42383 3556 42800 3584
rect 42383 3553 42395 3556
rect 42337 3547 42395 3553
rect 42794 3544 42800 3556
rect 42852 3544 42858 3596
rect 42904 3593 42932 3624
rect 45554 3612 45560 3624
rect 45612 3612 45618 3664
rect 45646 3612 45652 3664
rect 45704 3652 45710 3664
rect 47489 3655 47547 3661
rect 47489 3652 47501 3655
rect 45704 3624 47501 3652
rect 45704 3612 45710 3624
rect 47489 3621 47501 3624
rect 47535 3621 47547 3655
rect 47489 3615 47547 3621
rect 42889 3587 42947 3593
rect 42889 3553 42901 3587
rect 42935 3553 42947 3587
rect 42889 3547 42947 3553
rect 45189 3587 45247 3593
rect 45189 3553 45201 3587
rect 45235 3584 45247 3587
rect 48041 3587 48099 3593
rect 48041 3584 48053 3587
rect 45235 3556 48053 3584
rect 45235 3553 45247 3556
rect 45189 3547 45247 3553
rect 48041 3553 48053 3556
rect 48087 3553 48099 3587
rect 48041 3547 48099 3553
rect 45005 3519 45063 3525
rect 45005 3485 45017 3519
rect 45051 3485 45063 3519
rect 45005 3479 45063 3485
rect 47949 3519 48007 3525
rect 47949 3485 47961 3519
rect 47995 3516 48007 3519
rect 48148 3516 48176 3692
rect 47995 3488 48176 3516
rect 47995 3485 48007 3488
rect 47949 3479 48007 3485
rect 30374 3408 30380 3460
rect 30432 3448 30438 3460
rect 31389 3451 31447 3457
rect 31389 3448 31401 3451
rect 30432 3420 31401 3448
rect 30432 3408 30438 3420
rect 31389 3417 31401 3420
rect 31435 3417 31447 3451
rect 31389 3411 31447 3417
rect 34885 3451 34943 3457
rect 34885 3417 34897 3451
rect 34931 3448 34943 3451
rect 35434 3448 35440 3460
rect 34931 3420 35440 3448
rect 34931 3417 34943 3420
rect 34885 3411 34943 3417
rect 35434 3408 35440 3420
rect 35492 3408 35498 3460
rect 40037 3451 40095 3457
rect 40037 3417 40049 3451
rect 40083 3448 40095 3451
rect 40586 3448 40592 3460
rect 40083 3420 40592 3448
rect 40083 3417 40095 3420
rect 40037 3411 40095 3417
rect 40586 3408 40592 3420
rect 40644 3408 40650 3460
rect 37734 3380 37740 3392
rect 29472 3352 37740 3380
rect 28077 3343 28135 3349
rect 37734 3340 37740 3352
rect 37792 3340 37798 3392
rect 45020 3380 45048 3479
rect 45186 3408 45192 3460
rect 45244 3448 45250 3460
rect 46845 3451 46903 3457
rect 46845 3448 46857 3451
rect 45244 3420 46857 3448
rect 45244 3408 45250 3420
rect 46845 3417 46857 3420
rect 46891 3417 46903 3451
rect 46845 3411 46903 3417
rect 47762 3380 47768 3392
rect 45020 3352 47768 3380
rect 47762 3340 47768 3352
rect 47820 3340 47826 3392
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 2774 3176 2780 3188
rect 1688 3148 2780 3176
rect 1688 3049 1716 3148
rect 2774 3136 2780 3148
rect 2832 3136 2838 3188
rect 16666 3176 16672 3188
rect 6840 3148 16672 3176
rect 1857 3111 1915 3117
rect 1857 3077 1869 3111
rect 1903 3108 1915 3111
rect 3142 3108 3148 3120
rect 1903 3080 3148 3108
rect 1903 3077 1915 3080
rect 1857 3071 1915 3077
rect 3142 3068 3148 3080
rect 3200 3068 3206 3120
rect 4157 3111 4215 3117
rect 4157 3077 4169 3111
rect 4203 3108 4215 3111
rect 4614 3108 4620 3120
rect 4203 3080 4620 3108
rect 4203 3077 4215 3080
rect 4157 3071 4215 3077
rect 4614 3068 4620 3080
rect 4672 3068 4678 3120
rect 6840 3049 6868 3148
rect 16666 3136 16672 3148
rect 16724 3136 16730 3188
rect 21358 3176 21364 3188
rect 16868 3148 21364 3176
rect 7009 3111 7067 3117
rect 7009 3077 7021 3111
rect 7055 3108 7067 3111
rect 9030 3108 9036 3120
rect 7055 3080 9036 3108
rect 7055 3077 7067 3080
rect 7009 3071 7067 3077
rect 9030 3068 9036 3080
rect 9088 3068 9094 3120
rect 10965 3111 11023 3117
rect 10965 3077 10977 3111
rect 11011 3108 11023 3111
rect 12342 3108 12348 3120
rect 11011 3080 12348 3108
rect 11011 3077 11023 3080
rect 10965 3071 11023 3077
rect 12342 3068 12348 3080
rect 12400 3068 12406 3120
rect 14461 3111 14519 3117
rect 14461 3108 14473 3111
rect 14292 3080 14473 3108
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3009 1731 3043
rect 1673 3003 1731 3009
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 14182 3000 14188 3052
rect 14240 3040 14246 3052
rect 14292 3040 14320 3080
rect 14461 3077 14473 3080
rect 14507 3077 14519 3111
rect 16868 3108 16896 3148
rect 21358 3136 21364 3148
rect 21416 3136 21422 3188
rect 26206 3148 35894 3176
rect 17494 3108 17500 3120
rect 14461 3071 14519 3077
rect 15672 3080 16896 3108
rect 16960 3080 17500 3108
rect 14240 3012 14320 3040
rect 14240 3000 14246 3012
rect 2682 2972 2688 2984
rect 2643 2944 2688 2972
rect 2682 2932 2688 2944
rect 2740 2932 2746 2984
rect 3973 2975 4031 2981
rect 3973 2941 3985 2975
rect 4019 2972 4031 2975
rect 4798 2972 4804 2984
rect 4019 2944 4804 2972
rect 4019 2941 4031 2944
rect 3973 2935 4031 2941
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 5353 2975 5411 2981
rect 5353 2972 5365 2975
rect 5276 2944 5365 2972
rect 5276 2916 5304 2944
rect 5353 2941 5365 2944
rect 5399 2941 5411 2975
rect 5353 2935 5411 2941
rect 8665 2975 8723 2981
rect 8665 2941 8677 2975
rect 8711 2941 8723 2975
rect 8665 2935 8723 2941
rect 9125 2975 9183 2981
rect 9125 2941 9137 2975
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 9309 2975 9367 2981
rect 9309 2941 9321 2975
rect 9355 2972 9367 2975
rect 11054 2972 11060 2984
rect 9355 2944 11060 2972
rect 9355 2941 9367 2944
rect 9309 2935 9367 2941
rect 5258 2864 5264 2916
rect 5316 2864 5322 2916
rect 8680 2836 8708 2935
rect 9140 2904 9168 2935
rect 11054 2932 11060 2944
rect 11112 2932 11118 2984
rect 11977 2975 12035 2981
rect 11977 2941 11989 2975
rect 12023 2941 12035 2975
rect 12158 2972 12164 2984
rect 12119 2944 12164 2972
rect 11977 2935 12035 2941
rect 11882 2904 11888 2916
rect 9140 2876 11888 2904
rect 11882 2864 11888 2876
rect 11940 2864 11946 2916
rect 11054 2836 11060 2848
rect 8680 2808 11060 2836
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11992 2836 12020 2935
rect 12158 2932 12164 2944
rect 12216 2932 12222 2984
rect 13817 2975 13875 2981
rect 13817 2941 13829 2975
rect 13863 2972 13875 2975
rect 13998 2972 14004 2984
rect 13863 2944 14004 2972
rect 13863 2941 13875 2944
rect 13817 2935 13875 2941
rect 13998 2932 14004 2944
rect 14056 2932 14062 2984
rect 14277 2975 14335 2981
rect 14277 2941 14289 2975
rect 14323 2972 14335 2975
rect 15194 2972 15200 2984
rect 14323 2944 15200 2972
rect 14323 2941 14335 2944
rect 14277 2935 14335 2941
rect 15194 2932 15200 2944
rect 15252 2932 15258 2984
rect 12066 2864 12072 2916
rect 12124 2904 12130 2916
rect 14182 2904 14188 2916
rect 12124 2876 14188 2904
rect 12124 2864 12130 2876
rect 14182 2864 14188 2876
rect 14240 2864 14246 2916
rect 14550 2864 14556 2916
rect 14608 2904 14614 2916
rect 15672 2904 15700 3080
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3040 16175 3043
rect 16960 3040 16988 3080
rect 17494 3068 17500 3080
rect 17552 3068 17558 3120
rect 18969 3111 19027 3117
rect 18969 3077 18981 3111
rect 19015 3108 19027 3111
rect 19426 3108 19432 3120
rect 19015 3080 19432 3108
rect 19015 3077 19027 3080
rect 18969 3071 19027 3077
rect 19426 3068 19432 3080
rect 19484 3068 19490 3120
rect 19613 3111 19671 3117
rect 19613 3077 19625 3111
rect 19659 3108 19671 3111
rect 21450 3108 21456 3120
rect 19659 3080 21456 3108
rect 19659 3077 19671 3080
rect 19613 3071 19671 3077
rect 21450 3068 21456 3080
rect 21508 3068 21514 3120
rect 22462 3108 22468 3120
rect 22423 3080 22468 3108
rect 22462 3068 22468 3080
rect 22520 3068 22526 3120
rect 24762 3108 24768 3120
rect 24723 3080 24768 3108
rect 24762 3068 24768 3080
rect 24820 3068 24826 3120
rect 17126 3040 17132 3052
rect 16163 3012 16988 3040
rect 17087 3012 17132 3040
rect 16163 3009 16175 3012
rect 16117 3003 16175 3009
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 22278 3040 22284 3052
rect 22239 3012 22284 3040
rect 22278 3000 22284 3012
rect 22336 3000 22342 3052
rect 17313 2975 17371 2981
rect 17313 2941 17325 2975
rect 17359 2972 17371 2975
rect 17954 2972 17960 2984
rect 17359 2944 17960 2972
rect 17359 2941 17371 2944
rect 17313 2935 17371 2941
rect 17954 2932 17960 2944
rect 18012 2932 18018 2984
rect 19429 2975 19487 2981
rect 19429 2941 19441 2975
rect 19475 2972 19487 2975
rect 20806 2972 20812 2984
rect 19475 2944 20812 2972
rect 19475 2941 19487 2944
rect 19429 2935 19487 2941
rect 20806 2932 20812 2944
rect 20864 2932 20870 2984
rect 21269 2975 21327 2981
rect 21269 2941 21281 2975
rect 21315 2972 21327 2975
rect 21910 2972 21916 2984
rect 21315 2944 21916 2972
rect 21315 2941 21327 2944
rect 21269 2935 21327 2941
rect 21910 2932 21916 2944
rect 21968 2932 21974 2984
rect 23934 2972 23940 2984
rect 23895 2944 23940 2972
rect 23934 2932 23940 2944
rect 23992 2932 23998 2984
rect 24581 2975 24639 2981
rect 24581 2941 24593 2975
rect 24627 2972 24639 2975
rect 25314 2972 25320 2984
rect 24627 2944 25320 2972
rect 24627 2941 24639 2944
rect 24581 2935 24639 2941
rect 25314 2932 25320 2944
rect 25372 2932 25378 2984
rect 25958 2972 25964 2984
rect 25919 2944 25964 2972
rect 25958 2932 25964 2944
rect 26016 2932 26022 2984
rect 26206 2904 26234 3148
rect 27154 3108 27160 3120
rect 27115 3080 27160 3108
rect 27154 3068 27160 3080
rect 27212 3068 27218 3120
rect 29454 3108 29460 3120
rect 29415 3080 29460 3108
rect 29454 3068 29460 3080
rect 29512 3068 29518 3120
rect 32309 3111 32367 3117
rect 32309 3077 32321 3111
rect 32355 3108 32367 3111
rect 32398 3108 32404 3120
rect 32355 3080 32404 3108
rect 32355 3077 32367 3080
rect 32309 3071 32367 3077
rect 32398 3068 32404 3080
rect 32456 3068 32462 3120
rect 34606 3108 34612 3120
rect 34567 3080 34612 3108
rect 34606 3068 34612 3080
rect 34664 3068 34670 3120
rect 26970 3040 26976 3052
rect 26931 3012 26976 3040
rect 26970 3000 26976 3012
rect 27028 3000 27034 3052
rect 28902 3000 28908 3052
rect 28960 3040 28966 3052
rect 29273 3043 29331 3049
rect 29273 3040 29285 3043
rect 28960 3012 29285 3040
rect 28960 3000 28966 3012
rect 29273 3009 29285 3012
rect 29319 3009 29331 3043
rect 29273 3003 29331 3009
rect 31754 3000 31760 3052
rect 31812 3040 31818 3052
rect 32125 3043 32183 3049
rect 32125 3040 32137 3043
rect 31812 3012 32137 3040
rect 31812 3000 31818 3012
rect 32125 3009 32137 3012
rect 32171 3009 32183 3043
rect 32125 3003 32183 3009
rect 33594 3000 33600 3052
rect 33652 3040 33658 3052
rect 34422 3040 34428 3052
rect 33652 3012 34100 3040
rect 34383 3012 34428 3040
rect 33652 3000 33658 3012
rect 27154 2932 27160 2984
rect 27212 2972 27218 2984
rect 27433 2975 27491 2981
rect 27433 2972 27445 2975
rect 27212 2944 27445 2972
rect 27212 2932 27218 2944
rect 27433 2941 27445 2944
rect 27479 2941 27491 2975
rect 27433 2935 27491 2941
rect 29733 2975 29791 2981
rect 29733 2941 29745 2975
rect 29779 2941 29791 2975
rect 29733 2935 29791 2941
rect 32585 2975 32643 2981
rect 32585 2941 32597 2975
rect 32631 2941 32643 2975
rect 34072 2972 34100 3012
rect 34422 3000 34428 3012
rect 34480 3000 34486 3052
rect 34885 2975 34943 2981
rect 34885 2972 34897 2975
rect 34072 2944 34897 2972
rect 32585 2935 32643 2941
rect 34885 2941 34897 2944
rect 34931 2941 34943 2975
rect 34885 2935 34943 2941
rect 14608 2876 15700 2904
rect 17052 2876 26234 2904
rect 14608 2864 14614 2876
rect 17052 2836 17080 2876
rect 11992 2808 17080 2836
rect 21358 2796 21364 2848
rect 21416 2836 21422 2848
rect 28350 2836 28356 2848
rect 21416 2808 28356 2836
rect 21416 2796 21422 2808
rect 28350 2796 28356 2808
rect 28408 2796 28414 2848
rect 28442 2796 28448 2848
rect 28500 2836 28506 2848
rect 29748 2836 29776 2935
rect 28500 2808 29776 2836
rect 28500 2796 28506 2808
rect 31018 2796 31024 2848
rect 31076 2836 31082 2848
rect 32600 2836 32628 2935
rect 31076 2808 32628 2836
rect 35866 2836 35894 3148
rect 44744 3148 47808 3176
rect 37458 3108 37464 3120
rect 37419 3080 37464 3108
rect 37458 3068 37464 3080
rect 37516 3068 37522 3120
rect 38654 3068 38660 3120
rect 38712 3108 38718 3120
rect 39761 3111 39819 3117
rect 39761 3108 39773 3111
rect 38712 3080 39773 3108
rect 38712 3068 38718 3080
rect 39761 3077 39773 3080
rect 39807 3077 39819 3111
rect 39761 3071 39819 3077
rect 42058 3068 42064 3120
rect 42116 3108 42122 3120
rect 42613 3111 42671 3117
rect 42613 3108 42625 3111
rect 42116 3080 42625 3108
rect 42116 3068 42122 3080
rect 42613 3077 42625 3080
rect 42659 3077 42671 3111
rect 42613 3071 42671 3077
rect 39574 3040 39580 3052
rect 39535 3012 39580 3040
rect 39574 3000 39580 3012
rect 39632 3000 39638 3052
rect 42242 3000 42248 3052
rect 42300 3040 42306 3052
rect 42429 3043 42487 3049
rect 42429 3040 42441 3043
rect 42300 3012 42441 3040
rect 42300 3000 42306 3012
rect 42429 3009 42441 3012
rect 42475 3009 42487 3043
rect 42429 3003 42487 3009
rect 37277 2975 37335 2981
rect 37277 2941 37289 2975
rect 37323 2972 37335 2975
rect 37642 2972 37648 2984
rect 37323 2944 37648 2972
rect 37323 2941 37335 2944
rect 37277 2935 37335 2941
rect 37642 2932 37648 2944
rect 37700 2932 37706 2984
rect 37737 2975 37795 2981
rect 37737 2941 37749 2975
rect 37783 2941 37795 2975
rect 37737 2935 37795 2941
rect 36170 2864 36176 2916
rect 36228 2904 36234 2916
rect 37752 2904 37780 2935
rect 38746 2932 38752 2984
rect 38804 2972 38810 2984
rect 40037 2975 40095 2981
rect 40037 2972 40049 2975
rect 38804 2944 40049 2972
rect 38804 2932 38810 2944
rect 40037 2941 40049 2944
rect 40083 2941 40095 2975
rect 40037 2935 40095 2941
rect 41322 2932 41328 2984
rect 41380 2972 41386 2984
rect 44744 2981 44772 3148
rect 44910 3108 44916 3120
rect 44871 3080 44916 3108
rect 44910 3068 44916 3080
rect 44968 3068 44974 3120
rect 47780 3049 47808 3148
rect 47765 3043 47823 3049
rect 47765 3009 47777 3043
rect 47811 3009 47823 3043
rect 47765 3003 47823 3009
rect 42889 2975 42947 2981
rect 41380 2932 41414 2972
rect 42889 2941 42901 2975
rect 42935 2941 42947 2975
rect 42889 2935 42947 2941
rect 44729 2975 44787 2981
rect 44729 2941 44741 2975
rect 44775 2941 44787 2975
rect 44729 2935 44787 2941
rect 45189 2975 45247 2981
rect 45189 2941 45201 2975
rect 45235 2941 45247 2975
rect 45189 2935 45247 2941
rect 36228 2876 37780 2904
rect 41386 2904 41414 2932
rect 42904 2904 42932 2935
rect 41386 2876 42932 2904
rect 36228 2864 36234 2876
rect 42978 2836 42984 2848
rect 35866 2808 42984 2836
rect 31076 2796 31082 2808
rect 42978 2796 42984 2808
rect 43036 2796 43042 2848
rect 43898 2796 43904 2848
rect 43956 2836 43962 2848
rect 45204 2836 45232 2935
rect 43956 2808 45232 2836
rect 43956 2796 43962 2808
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 4614 2592 4620 2644
rect 4672 2592 4678 2644
rect 47762 2632 47768 2644
rect 47723 2604 47768 2632
rect 47762 2592 47768 2604
rect 47820 2592 47826 2644
rect 4632 2564 4660 2592
rect 10226 2564 10232 2576
rect 4172 2536 4660 2564
rect 8956 2536 10232 2564
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2456 1458 2508
rect 1581 2499 1639 2505
rect 1581 2465 1593 2499
rect 1627 2496 1639 2499
rect 1670 2496 1676 2508
rect 1627 2468 1676 2496
rect 1627 2465 1639 2468
rect 1581 2459 1639 2465
rect 1670 2456 1676 2468
rect 1728 2456 1734 2508
rect 2038 2496 2044 2508
rect 1999 2468 2044 2496
rect 2038 2456 2044 2468
rect 2096 2456 2102 2508
rect 3418 2456 3424 2508
rect 3476 2496 3482 2508
rect 4172 2505 4200 2536
rect 3973 2499 4031 2505
rect 3973 2496 3985 2499
rect 3476 2468 3985 2496
rect 3476 2456 3482 2468
rect 3973 2465 3985 2468
rect 4019 2465 4031 2499
rect 3973 2459 4031 2465
rect 4157 2499 4215 2505
rect 4157 2465 4169 2499
rect 4203 2465 4215 2499
rect 4614 2496 4620 2508
rect 4575 2468 4620 2496
rect 4157 2459 4215 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 6546 2496 6552 2508
rect 6507 2468 6552 2496
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 7742 2496 7748 2508
rect 7703 2468 7748 2496
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 8956 2505 8984 2536
rect 10226 2524 10232 2536
rect 10284 2524 10290 2576
rect 28810 2564 28816 2576
rect 16546 2536 26234 2564
rect 8941 2499 8999 2505
rect 8941 2465 8953 2499
rect 8987 2465 8999 2499
rect 8941 2459 8999 2465
rect 9122 2456 9128 2508
rect 9180 2496 9186 2508
rect 9401 2499 9459 2505
rect 9401 2496 9413 2499
rect 9180 2468 9413 2496
rect 9180 2456 9186 2468
rect 9401 2465 9413 2468
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 11609 2499 11667 2505
rect 11609 2465 11621 2499
rect 11655 2496 11667 2499
rect 16546 2496 16574 2536
rect 11655 2468 16574 2496
rect 11655 2465 11667 2468
rect 11609 2459 11667 2465
rect 16758 2456 16764 2508
rect 16816 2496 16822 2508
rect 16853 2499 16911 2505
rect 16853 2496 16865 2499
rect 16816 2468 16865 2496
rect 16816 2456 16822 2468
rect 16853 2465 16865 2468
rect 16899 2465 16911 2499
rect 17034 2496 17040 2508
rect 16995 2468 17040 2496
rect 16853 2459 16911 2465
rect 17034 2456 17040 2468
rect 17092 2456 17098 2508
rect 19334 2456 19340 2508
rect 19392 2496 19398 2508
rect 19429 2499 19487 2505
rect 19429 2496 19441 2499
rect 19392 2468 19441 2496
rect 19392 2456 19398 2468
rect 19429 2465 19441 2468
rect 19475 2465 19487 2499
rect 19429 2459 19487 2465
rect 19613 2499 19671 2505
rect 19613 2465 19625 2499
rect 19659 2496 19671 2499
rect 20346 2496 20352 2508
rect 19659 2468 20352 2496
rect 19659 2465 19671 2468
rect 19613 2459 19671 2465
rect 20346 2456 20352 2468
rect 20404 2456 20410 2508
rect 22002 2496 22008 2508
rect 21963 2468 22008 2496
rect 22002 2456 22008 2468
rect 22060 2456 22066 2508
rect 22189 2499 22247 2505
rect 22189 2465 22201 2499
rect 22235 2496 22247 2499
rect 23106 2496 23112 2508
rect 22235 2468 23112 2496
rect 22235 2465 22247 2468
rect 22189 2459 22247 2465
rect 23106 2456 23112 2468
rect 23164 2456 23170 2508
rect 23382 2456 23388 2508
rect 23440 2496 23446 2508
rect 23477 2499 23535 2505
rect 23477 2496 23489 2499
rect 23440 2468 23489 2496
rect 23440 2456 23446 2468
rect 23477 2465 23489 2468
rect 23523 2465 23535 2499
rect 24578 2496 24584 2508
rect 24539 2468 24584 2496
rect 23477 2459 23535 2465
rect 24578 2456 24584 2468
rect 24636 2456 24642 2508
rect 24765 2499 24823 2505
rect 24765 2465 24777 2499
rect 24811 2496 24823 2499
rect 25038 2496 25044 2508
rect 24811 2468 25044 2496
rect 24811 2465 24823 2468
rect 24765 2459 24823 2465
rect 25038 2456 25044 2468
rect 25096 2456 25102 2508
rect 25222 2496 25228 2508
rect 25183 2468 25228 2496
rect 25222 2456 25228 2468
rect 25280 2456 25286 2508
rect 13814 2428 13820 2440
rect 13004 2400 13820 2428
rect 6454 2320 6460 2372
rect 6512 2360 6518 2372
rect 6733 2363 6791 2369
rect 6733 2360 6745 2363
rect 6512 2332 6745 2360
rect 6512 2320 6518 2332
rect 6733 2329 6745 2332
rect 6779 2329 6791 2363
rect 6733 2323 6791 2329
rect 8846 2320 8852 2372
rect 8904 2360 8910 2372
rect 9125 2363 9183 2369
rect 9125 2360 9137 2363
rect 8904 2332 9137 2360
rect 8904 2320 8910 2332
rect 9125 2329 9137 2332
rect 9171 2329 9183 2363
rect 9125 2323 9183 2329
rect 11793 2363 11851 2369
rect 11793 2329 11805 2363
rect 11839 2360 11851 2363
rect 13004 2360 13032 2400
rect 13814 2388 13820 2400
rect 13872 2388 13878 2440
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 14148 2400 14289 2428
rect 14148 2388 14154 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 11839 2332 13032 2360
rect 13449 2363 13507 2369
rect 11839 2329 11851 2332
rect 11793 2323 11851 2329
rect 13449 2329 13461 2363
rect 13495 2360 13507 2363
rect 14461 2363 14519 2369
rect 13495 2332 14320 2360
rect 13495 2329 13507 2332
rect 13449 2323 13507 2329
rect 14292 2304 14320 2332
rect 14461 2329 14473 2363
rect 14507 2360 14519 2363
rect 15378 2360 15384 2372
rect 14507 2332 15384 2360
rect 14507 2329 14519 2332
rect 14461 2323 14519 2329
rect 15378 2320 15384 2332
rect 15436 2320 15442 2372
rect 16117 2363 16175 2369
rect 16117 2329 16129 2363
rect 16163 2360 16175 2363
rect 16850 2360 16856 2372
rect 16163 2332 16856 2360
rect 16163 2329 16175 2332
rect 16117 2323 16175 2329
rect 16850 2320 16856 2332
rect 16908 2320 16914 2372
rect 18693 2363 18751 2369
rect 18693 2329 18705 2363
rect 18739 2360 18751 2363
rect 18782 2360 18788 2372
rect 18739 2332 18788 2360
rect 18739 2329 18751 2332
rect 18693 2323 18751 2329
rect 18782 2320 18788 2332
rect 18840 2320 18846 2372
rect 21269 2363 21327 2369
rect 21269 2329 21281 2363
rect 21315 2360 21327 2363
rect 21358 2360 21364 2372
rect 21315 2332 21364 2360
rect 21315 2329 21327 2332
rect 21269 2323 21327 2329
rect 21358 2320 21364 2332
rect 21416 2320 21422 2372
rect 14274 2252 14280 2304
rect 14332 2252 14338 2304
rect 26206 2292 26234 2536
rect 26988 2536 28816 2564
rect 26988 2505 27016 2536
rect 28810 2524 28816 2536
rect 28868 2524 28874 2576
rect 29730 2524 29736 2576
rect 29788 2564 29794 2576
rect 29788 2536 30972 2564
rect 29788 2524 29794 2536
rect 26973 2499 27031 2505
rect 26973 2465 26985 2499
rect 27019 2465 27031 2499
rect 26973 2459 27031 2465
rect 27157 2499 27215 2505
rect 27157 2465 27169 2499
rect 27203 2496 27215 2499
rect 27614 2496 27620 2508
rect 27203 2468 27620 2496
rect 27203 2465 27215 2468
rect 27157 2459 27215 2465
rect 27614 2456 27620 2468
rect 27672 2456 27678 2508
rect 27798 2496 27804 2508
rect 27759 2468 27804 2496
rect 27798 2456 27804 2468
rect 27856 2456 27862 2508
rect 29549 2499 29607 2505
rect 29549 2465 29561 2499
rect 29595 2496 29607 2499
rect 30742 2496 30748 2508
rect 29595 2468 30748 2496
rect 29595 2465 29607 2468
rect 29549 2459 29607 2465
rect 30742 2456 30748 2468
rect 30800 2456 30806 2508
rect 30944 2505 30972 2536
rect 32214 2524 32220 2576
rect 32272 2564 32278 2576
rect 32272 2536 32352 2564
rect 32272 2524 32278 2536
rect 30929 2499 30987 2505
rect 30929 2465 30941 2499
rect 30975 2465 30987 2499
rect 30929 2459 30987 2465
rect 31938 2456 31944 2508
rect 31996 2496 32002 2508
rect 32324 2505 32352 2536
rect 37550 2524 37556 2576
rect 37608 2564 37614 2576
rect 37608 2536 38424 2564
rect 37608 2524 37614 2536
rect 32125 2499 32183 2505
rect 32125 2496 32137 2499
rect 31996 2468 32137 2496
rect 31996 2456 32002 2468
rect 32125 2465 32137 2468
rect 32171 2465 32183 2499
rect 32125 2459 32183 2465
rect 32309 2499 32367 2505
rect 32309 2465 32321 2499
rect 32355 2465 32367 2499
rect 32309 2459 32367 2465
rect 32398 2456 32404 2508
rect 32456 2496 32462 2508
rect 32585 2499 32643 2505
rect 32585 2496 32597 2499
rect 32456 2468 32597 2496
rect 32456 2456 32462 2468
rect 32585 2465 32597 2468
rect 32631 2465 32643 2499
rect 32585 2459 32643 2465
rect 34238 2456 34244 2508
rect 34296 2496 34302 2508
rect 35161 2499 35219 2505
rect 35161 2496 35173 2499
rect 34296 2468 35173 2496
rect 34296 2456 34302 2468
rect 35161 2465 35173 2468
rect 35207 2465 35219 2499
rect 37274 2496 37280 2508
rect 37235 2468 37280 2496
rect 35161 2459 35219 2465
rect 37274 2456 37280 2468
rect 37332 2456 37338 2508
rect 37461 2499 37519 2505
rect 37461 2465 37473 2499
rect 37507 2496 37519 2499
rect 38286 2496 38292 2508
rect 37507 2468 38292 2496
rect 37507 2465 37519 2468
rect 37461 2459 37519 2465
rect 38286 2456 38292 2468
rect 38344 2456 38350 2508
rect 38396 2505 38424 2536
rect 39482 2524 39488 2576
rect 39540 2564 39546 2576
rect 43530 2564 43536 2576
rect 39540 2536 40356 2564
rect 39540 2524 39546 2536
rect 38381 2499 38439 2505
rect 38381 2465 38393 2499
rect 38427 2465 38439 2499
rect 38381 2459 38439 2465
rect 39390 2456 39396 2508
rect 39448 2496 39454 2508
rect 39853 2499 39911 2505
rect 39853 2496 39865 2499
rect 39448 2468 39865 2496
rect 39448 2456 39454 2468
rect 39853 2465 39865 2468
rect 39899 2465 39911 2499
rect 40034 2496 40040 2508
rect 39995 2468 40040 2496
rect 39853 2459 39911 2465
rect 40034 2456 40040 2468
rect 40092 2456 40098 2508
rect 40328 2505 40356 2536
rect 42444 2536 43536 2564
rect 42444 2505 42472 2536
rect 43530 2524 43536 2536
rect 43588 2524 43594 2576
rect 44542 2524 44548 2576
rect 44600 2564 44606 2576
rect 44600 2536 45692 2564
rect 44600 2524 44606 2536
rect 40313 2499 40371 2505
rect 40313 2465 40325 2499
rect 40359 2465 40371 2499
rect 40313 2459 40371 2465
rect 42429 2499 42487 2505
rect 42429 2465 42441 2499
rect 42475 2465 42487 2499
rect 42610 2496 42616 2508
rect 42571 2468 42616 2496
rect 42429 2459 42487 2465
rect 42610 2456 42616 2468
rect 42668 2456 42674 2508
rect 42702 2456 42708 2508
rect 42760 2496 42766 2508
rect 42889 2499 42947 2505
rect 42889 2496 42901 2499
rect 42760 2468 42901 2496
rect 42760 2456 42766 2468
rect 42889 2465 42901 2468
rect 42935 2465 42947 2499
rect 42889 2459 42947 2465
rect 45005 2499 45063 2505
rect 45005 2465 45017 2499
rect 45051 2496 45063 2499
rect 45554 2496 45560 2508
rect 45051 2468 45560 2496
rect 45051 2465 45063 2468
rect 45005 2459 45063 2465
rect 45554 2456 45560 2468
rect 45612 2456 45618 2508
rect 45664 2505 45692 2536
rect 45649 2499 45707 2505
rect 45649 2465 45661 2499
rect 45695 2465 45707 2499
rect 45649 2459 45707 2465
rect 34698 2428 34704 2440
rect 34659 2400 34704 2428
rect 34698 2388 34704 2400
rect 34756 2388 34762 2440
rect 29086 2320 29092 2372
rect 29144 2360 29150 2372
rect 29733 2363 29791 2369
rect 29733 2360 29745 2363
rect 29144 2332 29745 2360
rect 29144 2320 29150 2332
rect 29733 2329 29745 2332
rect 29779 2329 29791 2363
rect 29733 2323 29791 2329
rect 34514 2320 34520 2372
rect 34572 2360 34578 2372
rect 34885 2363 34943 2369
rect 34885 2360 34897 2363
rect 34572 2332 34897 2360
rect 34572 2320 34578 2332
rect 34885 2329 34897 2332
rect 34931 2329 34943 2363
rect 34885 2323 34943 2329
rect 44450 2320 44456 2372
rect 44508 2360 44514 2372
rect 45189 2363 45247 2369
rect 45189 2360 45201 2363
rect 44508 2332 45201 2360
rect 44508 2320 44514 2332
rect 45189 2329 45201 2332
rect 45235 2329 45247 2363
rect 45189 2323 45247 2329
rect 38470 2292 38476 2304
rect 26206 2264 38476 2292
rect 38470 2252 38476 2264
rect 38528 2252 38534 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 13998 1504 14004 1556
rect 14056 1544 14062 1556
rect 14918 1544 14924 1556
rect 14056 1516 14924 1544
rect 14056 1504 14062 1516
rect 14918 1504 14924 1516
rect 14976 1504 14982 1556
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 2228 47132 2280 47184
rect 34888 47132 34940 47184
rect 1768 46996 1820 47048
rect 5264 47039 5316 47048
rect 5264 47005 5273 47039
rect 5273 47005 5307 47039
rect 5307 47005 5316 47039
rect 5264 46996 5316 47005
rect 21824 47039 21876 47048
rect 21824 47005 21833 47039
rect 21833 47005 21867 47039
rect 21867 47005 21876 47039
rect 21824 46996 21876 47005
rect 24952 46996 25004 47048
rect 28264 46996 28316 47048
rect 31760 46996 31812 47048
rect 34796 46996 34848 47048
rect 38200 46996 38252 47048
rect 44824 46996 44876 47048
rect 48136 46996 48188 47048
rect 8208 46928 8260 46980
rect 22008 46903 22060 46912
rect 22008 46869 22017 46903
rect 22017 46869 22051 46903
rect 22051 46869 22060 46903
rect 22008 46860 22060 46869
rect 25228 46903 25280 46912
rect 25228 46869 25237 46903
rect 25237 46869 25271 46903
rect 25271 46869 25280 46903
rect 25228 46860 25280 46869
rect 28540 46903 28592 46912
rect 28540 46869 28549 46903
rect 28549 46869 28583 46903
rect 28583 46869 28592 46903
rect 28540 46860 28592 46869
rect 32312 46903 32364 46912
rect 32312 46869 32321 46903
rect 32321 46869 32355 46903
rect 32355 46869 32364 46903
rect 32312 46860 32364 46869
rect 38476 46903 38528 46912
rect 38476 46869 38485 46903
rect 38485 46869 38519 46903
rect 38519 46869 38528 46903
rect 38476 46860 38528 46869
rect 41512 46860 41564 46912
rect 47952 46971 48004 46980
rect 47952 46937 47961 46971
rect 47961 46937 47995 46971
rect 47995 46937 48004 46971
rect 47952 46928 48004 46937
rect 42984 46903 43036 46912
rect 42984 46869 42993 46903
rect 42993 46869 43027 46903
rect 43027 46869 43036 46903
rect 42984 46860 43036 46869
rect 45560 46903 45612 46912
rect 45560 46869 45569 46903
rect 45569 46869 45603 46903
rect 45603 46869 45612 46903
rect 45560 46860 45612 46869
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 10324 8959 10376 8968
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 12532 8959 12584 8968
rect 10324 8916 10376 8925
rect 12532 8925 12541 8959
rect 12541 8925 12575 8959
rect 12575 8925 12584 8959
rect 12532 8916 12584 8925
rect 10416 8823 10468 8832
rect 10416 8789 10425 8823
rect 10425 8789 10459 8823
rect 10459 8789 10468 8823
rect 10416 8780 10468 8789
rect 11888 8780 11940 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 10968 8440 11020 8492
rect 47584 8440 47636 8492
rect 9588 8372 9640 8424
rect 1584 8304 1636 8356
rect 7748 8347 7800 8356
rect 7748 8313 7757 8347
rect 7757 8313 7791 8347
rect 7791 8313 7800 8347
rect 7748 8304 7800 8313
rect 8852 8304 8904 8356
rect 9036 8304 9088 8356
rect 9312 8304 9364 8356
rect 45376 8304 45428 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 8484 8032 8536 8084
rect 1400 7896 1452 7948
rect 10324 7896 10376 7948
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 6092 7871 6144 7880
rect 6092 7837 6101 7871
rect 6101 7837 6135 7871
rect 6135 7837 6144 7871
rect 6092 7828 6144 7837
rect 8208 7871 8260 7880
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 9588 7828 9640 7880
rect 10968 7871 11020 7880
rect 7196 7760 7248 7812
rect 7656 7760 7708 7812
rect 8944 7760 8996 7812
rect 10232 7760 10284 7812
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 47124 7871 47176 7880
rect 47124 7837 47133 7871
rect 47133 7837 47167 7871
rect 47167 7837 47176 7871
rect 47124 7828 47176 7837
rect 47584 7871 47636 7880
rect 47584 7837 47593 7871
rect 47593 7837 47627 7871
rect 47627 7837 47636 7871
rect 47584 7828 47636 7837
rect 47952 7760 48004 7812
rect 5172 7692 5224 7744
rect 7104 7735 7156 7744
rect 7104 7701 7113 7735
rect 7113 7701 7147 7735
rect 7147 7701 7156 7735
rect 7104 7692 7156 7701
rect 9220 7692 9272 7744
rect 11060 7735 11112 7744
rect 11060 7701 11069 7735
rect 11069 7701 11103 7735
rect 11103 7701 11112 7735
rect 11060 7692 11112 7701
rect 47676 7735 47728 7744
rect 47676 7701 47685 7735
rect 47685 7701 47719 7735
rect 47719 7701 47728 7735
rect 47676 7692 47728 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 5540 7352 5592 7404
rect 6092 7352 6144 7404
rect 6644 7352 6696 7404
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 8484 7420 8536 7472
rect 10416 7420 10468 7472
rect 10968 7352 11020 7404
rect 12440 7352 12492 7404
rect 47584 7395 47636 7404
rect 47584 7361 47593 7395
rect 47593 7361 47627 7395
rect 47627 7361 47636 7395
rect 47584 7352 47636 7361
rect 9496 7284 9548 7336
rect 45284 7284 45336 7336
rect 6368 7216 6420 7268
rect 11152 7216 11204 7268
rect 45468 7216 45520 7268
rect 1768 7148 1820 7200
rect 2780 7148 2832 7200
rect 5080 7191 5132 7200
rect 5080 7157 5089 7191
rect 5089 7157 5123 7191
rect 5123 7157 5132 7191
rect 5080 7148 5132 7157
rect 6460 7148 6512 7200
rect 7288 7191 7340 7200
rect 7288 7157 7297 7191
rect 7297 7157 7331 7191
rect 7331 7157 7340 7191
rect 7288 7148 7340 7157
rect 9864 7148 9916 7200
rect 11428 7148 11480 7200
rect 46388 7191 46440 7200
rect 46388 7157 46397 7191
rect 46397 7157 46431 7191
rect 46431 7157 46440 7191
rect 46388 7148 46440 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 5080 6944 5132 6996
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 3332 6740 3384 6792
rect 5540 6808 5592 6860
rect 5816 6808 5868 6860
rect 9496 6808 9548 6860
rect 10232 6808 10284 6860
rect 47124 6808 47176 6860
rect 4804 6740 4856 6792
rect 8944 6783 8996 6792
rect 4620 6672 4672 6724
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 9404 6740 9456 6792
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 12532 6740 12584 6792
rect 5724 6672 5776 6724
rect 7104 6672 7156 6724
rect 7564 6715 7616 6724
rect 7564 6681 7573 6715
rect 7573 6681 7607 6715
rect 7607 6681 7616 6715
rect 7564 6672 7616 6681
rect 10600 6715 10652 6724
rect 10600 6681 10609 6715
rect 10609 6681 10643 6715
rect 10643 6681 10652 6715
rect 10600 6672 10652 6681
rect 11888 6672 11940 6724
rect 47676 6672 47728 6724
rect 49056 6672 49108 6724
rect 2044 6647 2096 6656
rect 2044 6613 2053 6647
rect 2053 6613 2087 6647
rect 2087 6613 2096 6647
rect 2044 6604 2096 6613
rect 3148 6647 3200 6656
rect 3148 6613 3157 6647
rect 3157 6613 3191 6647
rect 3191 6613 3200 6647
rect 3148 6604 3200 6613
rect 4712 6604 4764 6656
rect 4988 6604 5040 6656
rect 5632 6604 5684 6656
rect 8024 6647 8076 6656
rect 8024 6613 8033 6647
rect 8033 6613 8067 6647
rect 8067 6613 8076 6647
rect 8024 6604 8076 6613
rect 9128 6604 9180 6656
rect 10324 6604 10376 6656
rect 13176 6647 13228 6656
rect 13176 6613 13185 6647
rect 13185 6613 13219 6647
rect 13219 6613 13228 6647
rect 13176 6604 13228 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 5080 6400 5132 6452
rect 8024 6400 8076 6452
rect 8116 6400 8168 6452
rect 9588 6400 9640 6452
rect 12440 6443 12492 6452
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 2596 6307 2648 6316
rect 1952 6264 2004 6273
rect 2596 6273 2605 6307
rect 2605 6273 2639 6307
rect 2639 6273 2648 6307
rect 2596 6264 2648 6273
rect 4068 6307 4120 6316
rect 4068 6273 4077 6307
rect 4077 6273 4111 6307
rect 4111 6273 4120 6307
rect 4068 6264 4120 6273
rect 4988 6264 5040 6316
rect 5264 6264 5316 6316
rect 9864 6332 9916 6384
rect 10232 6332 10284 6384
rect 12440 6409 12449 6443
rect 12449 6409 12483 6443
rect 12483 6409 12492 6443
rect 12440 6400 12492 6409
rect 1676 6060 1728 6112
rect 3608 6128 3660 6180
rect 4988 6128 5040 6180
rect 5724 6264 5776 6316
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 7748 6264 7800 6316
rect 8944 6264 8996 6316
rect 9496 6264 9548 6316
rect 9680 6307 9732 6316
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 10324 6307 10376 6316
rect 9680 6264 9732 6273
rect 10324 6273 10333 6307
rect 10333 6273 10367 6307
rect 10367 6273 10376 6307
rect 10324 6264 10376 6273
rect 12348 6307 12400 6316
rect 12348 6273 12357 6307
rect 12357 6273 12391 6307
rect 12391 6273 12400 6307
rect 12348 6264 12400 6273
rect 14372 6307 14424 6316
rect 14372 6273 14381 6307
rect 14381 6273 14415 6307
rect 14415 6273 14424 6307
rect 14372 6264 14424 6273
rect 46388 6332 46440 6384
rect 6644 6239 6696 6248
rect 6644 6205 6653 6239
rect 6653 6205 6687 6239
rect 6687 6205 6696 6239
rect 6644 6196 6696 6205
rect 6736 6196 6788 6248
rect 3424 6103 3476 6112
rect 3424 6069 3433 6103
rect 3433 6069 3467 6103
rect 3467 6069 3476 6103
rect 3424 6060 3476 6069
rect 3976 6060 4028 6112
rect 4896 6060 4948 6112
rect 7104 6060 7156 6112
rect 8668 6103 8720 6112
rect 8668 6069 8677 6103
rect 8677 6069 8711 6103
rect 8711 6069 8720 6103
rect 8668 6060 8720 6069
rect 9772 6196 9824 6248
rect 9404 6171 9456 6180
rect 9404 6137 9413 6171
rect 9413 6137 9447 6171
rect 9447 6137 9456 6171
rect 9404 6128 9456 6137
rect 10600 6196 10652 6248
rect 45376 6239 45428 6248
rect 45376 6205 45385 6239
rect 45385 6205 45419 6239
rect 45419 6205 45428 6239
rect 45376 6196 45428 6205
rect 48412 6196 48464 6248
rect 11796 6128 11848 6180
rect 13452 6128 13504 6180
rect 12440 6060 12492 6112
rect 13820 6103 13872 6112
rect 13820 6069 13829 6103
rect 13829 6069 13863 6103
rect 13863 6069 13872 6103
rect 13820 6060 13872 6069
rect 46296 6060 46348 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 6276 5856 6328 5908
rect 10232 5856 10284 5908
rect 11796 5899 11848 5908
rect 11796 5865 11805 5899
rect 11805 5865 11839 5899
rect 11839 5865 11848 5899
rect 11796 5856 11848 5865
rect 12440 5899 12492 5908
rect 12440 5865 12449 5899
rect 12449 5865 12483 5899
rect 12483 5865 12492 5899
rect 12440 5856 12492 5865
rect 8392 5788 8444 5840
rect 3240 5720 3292 5772
rect 3332 5652 3384 5704
rect 3700 5652 3752 5704
rect 4436 5695 4488 5704
rect 4436 5661 4445 5695
rect 4445 5661 4479 5695
rect 4479 5661 4488 5695
rect 4436 5652 4488 5661
rect 7288 5720 7340 5772
rect 7564 5720 7616 5772
rect 9680 5720 9732 5772
rect 10508 5720 10560 5772
rect 10692 5763 10744 5772
rect 10692 5729 10701 5763
rect 10701 5729 10735 5763
rect 10735 5729 10744 5763
rect 10692 5720 10744 5729
rect 11796 5720 11848 5772
rect 6368 5652 6420 5704
rect 8668 5652 8720 5704
rect 9496 5652 9548 5704
rect 9588 5652 9640 5704
rect 12348 5788 12400 5840
rect 13912 5788 13964 5840
rect 12440 5720 12492 5772
rect 31852 5720 31904 5772
rect 45836 5720 45888 5772
rect 46296 5763 46348 5772
rect 46296 5729 46305 5763
rect 46305 5729 46339 5763
rect 46339 5729 46348 5763
rect 46296 5720 46348 5729
rect 47124 5763 47176 5772
rect 47124 5729 47133 5763
rect 47133 5729 47167 5763
rect 47167 5729 47176 5763
rect 47124 5720 47176 5729
rect 14372 5652 14424 5704
rect 14924 5695 14976 5704
rect 14924 5661 14933 5695
rect 14933 5661 14967 5695
rect 14967 5661 14976 5695
rect 14924 5652 14976 5661
rect 31944 5652 31996 5704
rect 32128 5652 32180 5704
rect 36360 5695 36412 5704
rect 36360 5661 36369 5695
rect 36369 5661 36403 5695
rect 36403 5661 36412 5695
rect 36360 5652 36412 5661
rect 37280 5652 37332 5704
rect 39580 5652 39632 5704
rect 40132 5652 40184 5704
rect 41604 5695 41656 5704
rect 41604 5661 41613 5695
rect 41613 5661 41647 5695
rect 41647 5661 41656 5695
rect 41604 5652 41656 5661
rect 45008 5695 45060 5704
rect 45008 5661 45017 5695
rect 45017 5661 45051 5695
rect 45051 5661 45060 5695
rect 45008 5652 45060 5661
rect 45652 5695 45704 5704
rect 45652 5661 45661 5695
rect 45661 5661 45695 5695
rect 45695 5661 45704 5695
rect 45652 5652 45704 5661
rect 4252 5584 4304 5636
rect 4620 5584 4672 5636
rect 3792 5516 3844 5568
rect 4160 5516 4212 5568
rect 12164 5584 12216 5636
rect 6184 5559 6236 5568
rect 6184 5525 6193 5559
rect 6193 5525 6227 5559
rect 6227 5525 6236 5559
rect 6184 5516 6236 5525
rect 6828 5516 6880 5568
rect 7196 5516 7248 5568
rect 10508 5516 10560 5568
rect 14464 5516 14516 5568
rect 44916 5516 44968 5568
rect 45192 5516 45244 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4160 5312 4212 5364
rect 6644 5312 6696 5364
rect 6828 5312 6880 5364
rect 7196 5355 7248 5364
rect 7196 5321 7205 5355
rect 7205 5321 7239 5355
rect 7239 5321 7248 5355
rect 7196 5312 7248 5321
rect 7564 5312 7616 5364
rect 10324 5312 10376 5364
rect 10508 5355 10560 5364
rect 10508 5321 10517 5355
rect 10517 5321 10551 5355
rect 10551 5321 10560 5355
rect 10692 5355 10744 5364
rect 10508 5312 10560 5321
rect 10692 5321 10701 5355
rect 10701 5321 10735 5355
rect 10735 5321 10744 5355
rect 10692 5312 10744 5321
rect 2596 5244 2648 5296
rect 2320 5176 2372 5228
rect 2688 5176 2740 5228
rect 3700 5176 3752 5228
rect 5080 5244 5132 5296
rect 7104 5287 7156 5296
rect 7104 5253 7113 5287
rect 7113 5253 7147 5287
rect 7147 5253 7156 5287
rect 7104 5244 7156 5253
rect 8392 5244 8444 5296
rect 9128 5244 9180 5296
rect 9588 5244 9640 5296
rect 11796 5287 11848 5296
rect 11796 5253 11805 5287
rect 11805 5253 11839 5287
rect 11839 5253 11848 5287
rect 11796 5244 11848 5253
rect 13176 5244 13228 5296
rect 5632 5219 5684 5228
rect 5632 5185 5641 5219
rect 5641 5185 5675 5219
rect 5675 5185 5684 5219
rect 5632 5176 5684 5185
rect 10232 5176 10284 5228
rect 16488 5176 16540 5228
rect 18420 5176 18472 5228
rect 21088 5176 21140 5228
rect 28540 5176 28592 5228
rect 31668 5176 31720 5228
rect 33416 5219 33468 5228
rect 33416 5185 33425 5219
rect 33425 5185 33459 5219
rect 33459 5185 33468 5219
rect 33416 5176 33468 5185
rect 35440 5176 35492 5228
rect 37924 5219 37976 5228
rect 37924 5185 37933 5219
rect 37933 5185 37967 5219
rect 37967 5185 37976 5219
rect 37924 5176 37976 5185
rect 42432 5219 42484 5228
rect 42432 5185 42441 5219
rect 42441 5185 42475 5219
rect 42475 5185 42484 5219
rect 42432 5176 42484 5185
rect 45008 5176 45060 5228
rect 45468 5244 45520 5296
rect 47584 5219 47636 5228
rect 2872 5108 2924 5160
rect 5540 5151 5592 5160
rect 5540 5117 5549 5151
rect 5549 5117 5583 5151
rect 5583 5117 5592 5151
rect 5540 5108 5592 5117
rect 6552 5108 6604 5160
rect 7196 5108 7248 5160
rect 8484 5108 8536 5160
rect 45376 5151 45428 5160
rect 45376 5117 45385 5151
rect 45385 5117 45419 5151
rect 45419 5117 45428 5151
rect 45376 5108 45428 5117
rect 45652 5108 45704 5160
rect 47584 5185 47593 5219
rect 47593 5185 47627 5219
rect 47627 5185 47636 5219
rect 47584 5176 47636 5185
rect 47676 5108 47728 5160
rect 3976 5040 4028 5092
rect 5816 5040 5868 5092
rect 3056 5015 3108 5024
rect 3056 4981 3065 5015
rect 3065 4981 3099 5015
rect 3099 4981 3108 5015
rect 3056 4972 3108 4981
rect 9496 4972 9548 5024
rect 14096 5040 14148 5092
rect 32404 5040 32456 5092
rect 34612 5040 34664 5092
rect 37648 5040 37700 5092
rect 14372 5015 14424 5024
rect 14372 4981 14381 5015
rect 14381 4981 14415 5015
rect 14415 4981 14424 5015
rect 14372 4972 14424 4981
rect 15200 4972 15252 5024
rect 15936 4972 15988 5024
rect 17408 5015 17460 5024
rect 17408 4981 17417 5015
rect 17417 4981 17451 5015
rect 17451 4981 17460 5015
rect 17408 4972 17460 4981
rect 17960 4972 18012 5024
rect 19156 5015 19208 5024
rect 19156 4981 19165 5015
rect 19165 4981 19199 5015
rect 19199 4981 19208 5015
rect 19156 4972 19208 4981
rect 19340 4972 19392 5024
rect 20352 5015 20404 5024
rect 20352 4981 20361 5015
rect 20361 4981 20395 5015
rect 20395 4981 20404 5015
rect 20352 4972 20404 4981
rect 20812 4972 20864 5024
rect 21456 4972 21508 5024
rect 22284 4972 22336 5024
rect 23848 4972 23900 5024
rect 24584 4972 24636 5024
rect 28448 5015 28500 5024
rect 28448 4981 28457 5015
rect 28457 4981 28491 5015
rect 28491 4981 28500 5015
rect 28448 4972 28500 4981
rect 29092 5015 29144 5024
rect 29092 4981 29101 5015
rect 29101 4981 29135 5015
rect 29135 4981 29144 5015
rect 29092 4972 29144 4981
rect 32036 4972 32088 5024
rect 32220 5015 32272 5024
rect 32220 4981 32229 5015
rect 32229 4981 32263 5015
rect 32263 4981 32272 5015
rect 32220 4972 32272 4981
rect 32312 4972 32364 5024
rect 34520 4972 34572 5024
rect 34704 4972 34756 5024
rect 35348 4972 35400 5024
rect 37372 5015 37424 5024
rect 37372 4981 37381 5015
rect 37381 4981 37415 5015
rect 37415 4981 37424 5015
rect 37372 4972 37424 4981
rect 37556 4972 37608 5024
rect 38660 5015 38712 5024
rect 38660 4981 38669 5015
rect 38669 4981 38703 5015
rect 38703 4981 38712 5015
rect 38660 4972 38712 4981
rect 39396 5015 39448 5024
rect 39396 4981 39405 5015
rect 39405 4981 39439 5015
rect 39439 4981 39448 5015
rect 39396 4972 39448 4981
rect 40224 4972 40276 5024
rect 40592 5015 40644 5024
rect 40592 4981 40601 5015
rect 40601 4981 40635 5015
rect 40635 4981 40644 5015
rect 40592 4972 40644 4981
rect 42064 4972 42116 5024
rect 42616 4972 42668 5024
rect 43260 5015 43312 5024
rect 43260 4981 43269 5015
rect 43269 4981 43303 5015
rect 43303 4981 43312 5015
rect 43260 4972 43312 4981
rect 43812 5015 43864 5024
rect 43812 4981 43821 5015
rect 43821 4981 43855 5015
rect 43855 4981 43864 5015
rect 43812 4972 43864 4981
rect 44456 5015 44508 5024
rect 44456 4981 44465 5015
rect 44465 4981 44499 5015
rect 44499 4981 44508 5015
rect 44456 4972 44508 4981
rect 46020 4972 46072 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 4068 4768 4120 4820
rect 31668 4768 31720 4820
rect 33416 4768 33468 4820
rect 45652 4768 45704 4820
rect 2872 4675 2924 4684
rect 2872 4641 2881 4675
rect 2881 4641 2915 4675
rect 2915 4641 2924 4675
rect 2872 4632 2924 4641
rect 2688 4564 2740 4616
rect 4896 4700 4948 4752
rect 3240 4632 3292 4684
rect 4252 4675 4304 4684
rect 4252 4641 4261 4675
rect 4261 4641 4295 4675
rect 4295 4641 4304 4675
rect 4252 4632 4304 4641
rect 5540 4632 5592 4684
rect 6184 4632 6236 4684
rect 6460 4675 6512 4684
rect 6460 4641 6469 4675
rect 6469 4641 6503 4675
rect 6503 4641 6512 4675
rect 6460 4632 6512 4641
rect 6920 4675 6972 4684
rect 6920 4641 6929 4675
rect 6929 4641 6963 4675
rect 6963 4641 6972 4675
rect 6920 4632 6972 4641
rect 10324 4700 10376 4752
rect 14924 4700 14976 4752
rect 24952 4700 25004 4752
rect 9220 4632 9272 4684
rect 9772 4675 9824 4684
rect 9772 4641 9781 4675
rect 9781 4641 9815 4675
rect 9815 4641 9824 4675
rect 9772 4632 9824 4641
rect 34796 4700 34848 4752
rect 28908 4632 28960 4684
rect 45836 4675 45888 4684
rect 15844 4564 15896 4616
rect 16120 4607 16172 4616
rect 16120 4573 16129 4607
rect 16129 4573 16163 4607
rect 16163 4573 16172 4607
rect 16120 4564 16172 4573
rect 16764 4607 16816 4616
rect 16764 4573 16773 4607
rect 16773 4573 16807 4607
rect 16807 4573 16816 4607
rect 16764 4564 16816 4573
rect 17132 4564 17184 4616
rect 18052 4607 18104 4616
rect 18052 4573 18061 4607
rect 18061 4573 18095 4607
rect 18095 4573 18104 4607
rect 18052 4564 18104 4573
rect 18420 4564 18472 4616
rect 20536 4607 20588 4616
rect 2872 4496 2924 4548
rect 3608 4496 3660 4548
rect 12440 4496 12492 4548
rect 13636 4496 13688 4548
rect 14648 4496 14700 4548
rect 19432 4496 19484 4548
rect 20536 4573 20545 4607
rect 20545 4573 20579 4607
rect 20579 4573 20588 4607
rect 20536 4564 20588 4573
rect 21916 4607 21968 4616
rect 21916 4573 21925 4607
rect 21925 4573 21959 4607
rect 21959 4573 21968 4607
rect 21916 4564 21968 4573
rect 21088 4496 21140 4548
rect 23296 4564 23348 4616
rect 25320 4564 25372 4616
rect 27620 4564 27672 4616
rect 28540 4607 28592 4616
rect 28540 4573 28549 4607
rect 28549 4573 28583 4607
rect 28583 4573 28592 4607
rect 28540 4564 28592 4573
rect 29736 4607 29788 4616
rect 29736 4573 29745 4607
rect 29745 4573 29779 4607
rect 29779 4573 29788 4607
rect 29736 4564 29788 4573
rect 30380 4607 30432 4616
rect 30380 4573 30389 4607
rect 30389 4573 30423 4607
rect 30423 4573 30432 4607
rect 30380 4564 30432 4573
rect 31760 4564 31812 4616
rect 34428 4564 34480 4616
rect 34796 4564 34848 4616
rect 35440 4564 35492 4616
rect 36176 4607 36228 4616
rect 36176 4573 36185 4607
rect 36185 4573 36219 4607
rect 36219 4573 36228 4607
rect 36176 4564 36228 4573
rect 23388 4496 23440 4548
rect 37924 4564 37976 4616
rect 39028 4607 39080 4616
rect 39028 4573 39037 4607
rect 39037 4573 39071 4607
rect 39071 4573 39080 4607
rect 39028 4564 39080 4573
rect 42248 4607 42300 4616
rect 42248 4573 42257 4607
rect 42257 4573 42291 4607
rect 42291 4573 42300 4607
rect 42248 4564 42300 4573
rect 42432 4564 42484 4616
rect 43536 4607 43588 4616
rect 43536 4573 43545 4607
rect 43545 4573 43579 4607
rect 43579 4573 43588 4607
rect 43536 4564 43588 4573
rect 45836 4641 45845 4675
rect 45845 4641 45879 4675
rect 45879 4641 45888 4675
rect 45836 4632 45888 4641
rect 46020 4675 46072 4684
rect 46020 4641 46029 4675
rect 46029 4641 46063 4675
rect 46063 4641 46072 4675
rect 46020 4632 46072 4641
rect 46480 4675 46532 4684
rect 46480 4641 46489 4675
rect 46489 4641 46523 4675
rect 46523 4641 46532 4675
rect 46480 4632 46532 4641
rect 2228 4428 2280 4480
rect 6460 4428 6512 4480
rect 15384 4471 15436 4480
rect 15384 4437 15393 4471
rect 15393 4437 15427 4471
rect 15427 4437 15436 4471
rect 15384 4428 15436 4437
rect 18696 4428 18748 4480
rect 22100 4428 22152 4480
rect 23112 4471 23164 4480
rect 23112 4437 23121 4471
rect 23121 4437 23155 4471
rect 23155 4437 23164 4471
rect 23112 4428 23164 4437
rect 24032 4428 24084 4480
rect 24768 4428 24820 4480
rect 25872 4428 25924 4480
rect 29460 4428 29512 4480
rect 35440 4471 35492 4480
rect 35440 4437 35449 4471
rect 35449 4437 35483 4471
rect 35483 4437 35492 4471
rect 35440 4428 35492 4437
rect 37464 4428 37516 4480
rect 45008 4496 45060 4548
rect 45376 4539 45428 4548
rect 45376 4505 45385 4539
rect 45385 4505 45419 4539
rect 45419 4505 45428 4539
rect 45376 4496 45428 4505
rect 37740 4428 37792 4480
rect 38292 4471 38344 4480
rect 38292 4437 38301 4471
rect 38301 4437 38335 4471
rect 38335 4437 38344 4471
rect 38292 4428 38344 4437
rect 40040 4428 40092 4480
rect 41512 4471 41564 4480
rect 41512 4437 41521 4471
rect 41521 4437 41555 4471
rect 41555 4437 41564 4471
rect 41512 4428 41564 4437
rect 42800 4471 42852 4480
rect 42800 4437 42809 4471
rect 42809 4437 42843 4471
rect 42843 4437 42852 4471
rect 42800 4428 42852 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2228 4224 2280 4276
rect 5540 4224 5592 4276
rect 20536 4224 20588 4276
rect 23296 4267 23348 4276
rect 2320 4156 2372 4208
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 756 3952 808 4004
rect 3792 4020 3844 4072
rect 7012 4063 7064 4072
rect 3332 3952 3384 4004
rect 4252 3952 4304 4004
rect 3976 3884 4028 3936
rect 7012 4029 7021 4063
rect 7021 4029 7055 4063
rect 7055 4029 7064 4063
rect 7012 4020 7064 4029
rect 7196 4020 7248 4072
rect 9312 4063 9364 4072
rect 7104 3952 7156 4004
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 11704 4020 11756 4072
rect 13912 4156 13964 4208
rect 14648 4156 14700 4208
rect 15844 4131 15896 4140
rect 15844 4097 15853 4131
rect 15853 4097 15887 4131
rect 15887 4097 15896 4131
rect 15844 4088 15896 4097
rect 16488 4088 16540 4140
rect 18420 4156 18472 4208
rect 18696 4199 18748 4208
rect 18696 4165 18705 4199
rect 18705 4165 18739 4199
rect 18739 4165 18748 4199
rect 18696 4156 18748 4165
rect 21088 4199 21140 4208
rect 21088 4165 21097 4199
rect 21097 4165 21131 4199
rect 21131 4165 21140 4199
rect 21088 4156 21140 4165
rect 18052 4088 18104 4140
rect 23296 4233 23305 4267
rect 23305 4233 23339 4267
rect 23339 4233 23348 4267
rect 23296 4224 23348 4233
rect 23388 4156 23440 4208
rect 24032 4199 24084 4208
rect 24032 4165 24041 4199
rect 24041 4165 24075 4199
rect 24075 4165 24084 4199
rect 24032 4156 24084 4165
rect 28448 4199 28500 4208
rect 28448 4165 28457 4199
rect 28457 4165 28491 4199
rect 28491 4165 28500 4199
rect 28448 4156 28500 4165
rect 32312 4199 32364 4208
rect 32312 4165 32321 4199
rect 32321 4165 32355 4199
rect 32355 4165 32364 4199
rect 32312 4156 32364 4165
rect 35348 4156 35400 4208
rect 37556 4199 37608 4208
rect 37556 4165 37565 4199
rect 37565 4165 37599 4199
rect 37599 4165 37608 4199
rect 37556 4156 37608 4165
rect 23848 4131 23900 4140
rect 13084 4063 13136 4072
rect 13084 4029 13093 4063
rect 13093 4029 13127 4063
rect 13127 4029 13136 4063
rect 13084 4020 13136 4029
rect 13268 4063 13320 4072
rect 13268 4029 13277 4063
rect 13277 4029 13311 4063
rect 13311 4029 13320 4063
rect 13268 4020 13320 4029
rect 13452 4063 13504 4072
rect 13452 4029 13461 4063
rect 13461 4029 13495 4063
rect 13495 4029 13504 4063
rect 13452 4020 13504 4029
rect 15568 4020 15620 4072
rect 20076 4063 20128 4072
rect 20076 4029 20085 4063
rect 20085 4029 20119 4063
rect 20119 4029 20128 4063
rect 20076 4020 20128 4029
rect 23848 4097 23857 4131
rect 23857 4097 23891 4131
rect 23891 4097 23900 4131
rect 23848 4088 23900 4097
rect 27620 4131 27672 4140
rect 27620 4097 27629 4131
rect 27629 4097 27663 4131
rect 27663 4097 27672 4131
rect 27620 4088 27672 4097
rect 31668 4088 31720 4140
rect 32128 4131 32180 4140
rect 32128 4097 32137 4131
rect 32137 4097 32171 4131
rect 32171 4097 32180 4131
rect 32128 4088 32180 4097
rect 43260 4156 43312 4208
rect 23296 4020 23348 4072
rect 24492 4063 24544 4072
rect 24492 4029 24501 4063
rect 24501 4029 24535 4063
rect 24535 4029 24544 4063
rect 24492 4020 24544 4029
rect 29736 4020 29788 4072
rect 32956 4063 33008 4072
rect 25228 3952 25280 4004
rect 26240 3952 26292 4004
rect 13084 3884 13136 3936
rect 16304 3884 16356 3936
rect 17040 3884 17092 3936
rect 19432 3884 19484 3936
rect 22008 3927 22060 3936
rect 22008 3893 22017 3927
rect 22017 3893 22051 3927
rect 22051 3893 22060 3927
rect 22008 3884 22060 3893
rect 22468 3884 22520 3936
rect 25688 3884 25740 3936
rect 26976 3884 27028 3936
rect 27620 3884 27672 3936
rect 29184 3952 29236 4004
rect 32956 4029 32965 4063
rect 32965 4029 32999 4063
rect 32999 4029 33008 4063
rect 32956 4020 33008 4029
rect 32496 3952 32548 4004
rect 36176 4020 36228 4072
rect 38108 4063 38160 4072
rect 35532 3952 35584 4004
rect 38108 4029 38117 4063
rect 38117 4029 38151 4063
rect 38151 4029 38160 4063
rect 38108 4020 38160 4029
rect 39028 3952 39080 4004
rect 41512 4020 41564 4072
rect 40132 3952 40184 4004
rect 40684 3952 40736 4004
rect 43812 4020 43864 4072
rect 45192 4063 45244 4072
rect 43260 3952 43312 4004
rect 45192 4029 45201 4063
rect 45201 4029 45235 4063
rect 45235 4029 45244 4063
rect 45192 4020 45244 4029
rect 45836 4063 45888 4072
rect 45836 4029 45845 4063
rect 45845 4029 45879 4063
rect 45879 4029 45888 4063
rect 45836 4020 45888 4029
rect 30748 3927 30800 3936
rect 30748 3893 30757 3927
rect 30757 3893 30791 3927
rect 30791 3893 30800 3927
rect 30748 3884 30800 3893
rect 31300 3927 31352 3936
rect 31300 3893 31309 3927
rect 31309 3893 31343 3927
rect 31343 3893 31352 3927
rect 31300 3884 31352 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 1860 3680 1912 3732
rect 13268 3680 13320 3732
rect 2872 3612 2924 3664
rect 1584 3544 1636 3596
rect 4988 3612 5040 3664
rect 5172 3544 5224 3596
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 9496 3612 9548 3664
rect 9588 3544 9640 3596
rect 10416 3587 10468 3596
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 14372 3544 14424 3596
rect 16120 3544 16172 3596
rect 17408 3544 17460 3596
rect 18144 3587 18196 3596
rect 18144 3553 18153 3587
rect 18153 3553 18187 3587
rect 18187 3553 18196 3587
rect 18144 3544 18196 3553
rect 19156 3544 19208 3596
rect 19432 3587 19484 3596
rect 19432 3553 19441 3587
rect 19441 3553 19475 3587
rect 19475 3553 19484 3587
rect 19432 3544 19484 3553
rect 20720 3587 20772 3596
rect 20720 3553 20729 3587
rect 20729 3553 20763 3587
rect 20763 3553 20772 3587
rect 20720 3544 20772 3553
rect 21916 3544 21968 3596
rect 24952 3612 25004 3664
rect 26240 3544 26292 3596
rect 26516 3587 26568 3596
rect 26516 3553 26525 3587
rect 26525 3553 26559 3587
rect 26559 3553 26568 3587
rect 26516 3544 26568 3553
rect 24952 3519 25004 3528
rect 24952 3485 24961 3519
rect 24961 3485 24995 3519
rect 24995 3485 25004 3519
rect 24952 3476 25004 3485
rect 25688 3519 25740 3528
rect 25688 3485 25697 3519
rect 25697 3485 25731 3519
rect 25731 3485 25740 3519
rect 25688 3476 25740 3485
rect 27712 3476 27764 3528
rect 28816 3519 28868 3528
rect 28816 3485 28825 3519
rect 28825 3485 28859 3519
rect 28859 3485 28868 3519
rect 28816 3476 28868 3485
rect 2044 3408 2096 3460
rect 6276 3408 6328 3460
rect 8484 3408 8536 3460
rect 11152 3408 11204 3460
rect 11428 3451 11480 3460
rect 11428 3417 11437 3451
rect 11437 3417 11471 3451
rect 11471 3417 11480 3451
rect 11428 3408 11480 3417
rect 12992 3408 13044 3460
rect 14464 3408 14516 3460
rect 16212 3408 16264 3460
rect 16304 3408 16356 3460
rect 19524 3408 19576 3460
rect 22100 3408 22152 3460
rect 22652 3408 22704 3460
rect 25872 3451 25924 3460
rect 25872 3417 25881 3451
rect 25881 3417 25915 3451
rect 25915 3417 25924 3451
rect 25872 3408 25924 3417
rect 14188 3340 14240 3392
rect 15936 3340 15988 3392
rect 16672 3340 16724 3392
rect 21732 3340 21784 3392
rect 25044 3383 25096 3392
rect 25044 3349 25053 3383
rect 25053 3349 25087 3383
rect 25087 3349 25096 3383
rect 25044 3340 25096 3349
rect 27160 3340 27212 3392
rect 30380 3612 30432 3664
rect 31668 3612 31720 3664
rect 31300 3544 31352 3596
rect 31852 3587 31904 3596
rect 31852 3553 31861 3587
rect 31861 3553 31895 3587
rect 31895 3553 31904 3587
rect 31852 3544 31904 3553
rect 32036 3587 32088 3596
rect 32036 3553 32045 3587
rect 32045 3553 32079 3587
rect 32079 3553 32088 3587
rect 32036 3544 32088 3553
rect 36820 3612 36872 3664
rect 34704 3587 34756 3596
rect 34704 3553 34713 3587
rect 34713 3553 34747 3587
rect 34747 3553 34756 3587
rect 34704 3544 34756 3553
rect 34888 3544 34940 3596
rect 36360 3544 36412 3596
rect 37372 3544 37424 3596
rect 40132 3612 40184 3664
rect 40224 3544 40276 3596
rect 41972 3612 42024 3664
rect 45376 3680 45428 3732
rect 41604 3544 41656 3596
rect 42800 3544 42852 3596
rect 45560 3612 45612 3664
rect 45652 3612 45704 3664
rect 30380 3408 30432 3460
rect 35440 3408 35492 3460
rect 40592 3408 40644 3460
rect 37740 3340 37792 3392
rect 45192 3408 45244 3460
rect 47768 3340 47820 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2780 3136 2832 3188
rect 3148 3068 3200 3120
rect 4620 3068 4672 3120
rect 16672 3136 16724 3188
rect 9036 3068 9088 3120
rect 12348 3068 12400 3120
rect 14188 3000 14240 3052
rect 21364 3136 21416 3188
rect 2688 2975 2740 2984
rect 2688 2941 2697 2975
rect 2697 2941 2731 2975
rect 2731 2941 2740 2975
rect 2688 2932 2740 2941
rect 4804 2932 4856 2984
rect 5264 2864 5316 2916
rect 11060 2932 11112 2984
rect 12164 2975 12216 2984
rect 11888 2864 11940 2916
rect 11060 2796 11112 2848
rect 12164 2941 12173 2975
rect 12173 2941 12207 2975
rect 12207 2941 12216 2975
rect 12164 2932 12216 2941
rect 14004 2932 14056 2984
rect 15200 2932 15252 2984
rect 12072 2864 12124 2916
rect 14188 2864 14240 2916
rect 14556 2864 14608 2916
rect 17500 3068 17552 3120
rect 19432 3068 19484 3120
rect 21456 3068 21508 3120
rect 22468 3111 22520 3120
rect 22468 3077 22477 3111
rect 22477 3077 22511 3111
rect 22511 3077 22520 3111
rect 22468 3068 22520 3077
rect 24768 3111 24820 3120
rect 24768 3077 24777 3111
rect 24777 3077 24811 3111
rect 24811 3077 24820 3111
rect 24768 3068 24820 3077
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 22284 3043 22336 3052
rect 22284 3009 22293 3043
rect 22293 3009 22327 3043
rect 22327 3009 22336 3043
rect 22284 3000 22336 3009
rect 17960 2932 18012 2984
rect 20812 2932 20864 2984
rect 21916 2932 21968 2984
rect 23940 2975 23992 2984
rect 23940 2941 23949 2975
rect 23949 2941 23983 2975
rect 23983 2941 23992 2975
rect 23940 2932 23992 2941
rect 25320 2932 25372 2984
rect 25964 2975 26016 2984
rect 25964 2941 25973 2975
rect 25973 2941 26007 2975
rect 26007 2941 26016 2975
rect 25964 2932 26016 2941
rect 27160 3111 27212 3120
rect 27160 3077 27169 3111
rect 27169 3077 27203 3111
rect 27203 3077 27212 3111
rect 27160 3068 27212 3077
rect 29460 3111 29512 3120
rect 29460 3077 29469 3111
rect 29469 3077 29503 3111
rect 29503 3077 29512 3111
rect 29460 3068 29512 3077
rect 32404 3068 32456 3120
rect 34612 3111 34664 3120
rect 34612 3077 34621 3111
rect 34621 3077 34655 3111
rect 34655 3077 34664 3111
rect 34612 3068 34664 3077
rect 26976 3043 27028 3052
rect 26976 3009 26985 3043
rect 26985 3009 27019 3043
rect 27019 3009 27028 3043
rect 26976 3000 27028 3009
rect 28908 3000 28960 3052
rect 31760 3000 31812 3052
rect 33600 3000 33652 3052
rect 34428 3043 34480 3052
rect 27160 2932 27212 2984
rect 34428 3009 34437 3043
rect 34437 3009 34471 3043
rect 34471 3009 34480 3043
rect 34428 3000 34480 3009
rect 21364 2796 21416 2848
rect 28356 2796 28408 2848
rect 28448 2796 28500 2848
rect 31024 2796 31076 2848
rect 37464 3111 37516 3120
rect 37464 3077 37473 3111
rect 37473 3077 37507 3111
rect 37507 3077 37516 3111
rect 37464 3068 37516 3077
rect 38660 3068 38712 3120
rect 42064 3068 42116 3120
rect 39580 3043 39632 3052
rect 39580 3009 39589 3043
rect 39589 3009 39623 3043
rect 39623 3009 39632 3043
rect 39580 3000 39632 3009
rect 42248 3000 42300 3052
rect 37648 2932 37700 2984
rect 36176 2864 36228 2916
rect 38752 2932 38804 2984
rect 41328 2932 41380 2984
rect 44916 3111 44968 3120
rect 44916 3077 44925 3111
rect 44925 3077 44959 3111
rect 44959 3077 44968 3111
rect 44916 3068 44968 3077
rect 42984 2796 43036 2848
rect 43904 2796 43956 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4620 2592 4672 2644
rect 47768 2635 47820 2644
rect 47768 2601 47777 2635
rect 47777 2601 47811 2635
rect 47811 2601 47820 2635
rect 47768 2592 47820 2601
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 1676 2456 1728 2508
rect 2044 2499 2096 2508
rect 2044 2465 2053 2499
rect 2053 2465 2087 2499
rect 2087 2465 2096 2499
rect 2044 2456 2096 2465
rect 3424 2456 3476 2508
rect 4620 2499 4672 2508
rect 4620 2465 4629 2499
rect 4629 2465 4663 2499
rect 4663 2465 4672 2499
rect 4620 2456 4672 2465
rect 6552 2499 6604 2508
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 7748 2499 7800 2508
rect 7748 2465 7757 2499
rect 7757 2465 7791 2499
rect 7791 2465 7800 2499
rect 7748 2456 7800 2465
rect 10232 2524 10284 2576
rect 9128 2456 9180 2508
rect 16764 2456 16816 2508
rect 17040 2499 17092 2508
rect 17040 2465 17049 2499
rect 17049 2465 17083 2499
rect 17083 2465 17092 2499
rect 17040 2456 17092 2465
rect 19340 2456 19392 2508
rect 20352 2456 20404 2508
rect 22008 2499 22060 2508
rect 22008 2465 22017 2499
rect 22017 2465 22051 2499
rect 22051 2465 22060 2499
rect 22008 2456 22060 2465
rect 23112 2456 23164 2508
rect 23388 2456 23440 2508
rect 24584 2499 24636 2508
rect 24584 2465 24593 2499
rect 24593 2465 24627 2499
rect 24627 2465 24636 2499
rect 24584 2456 24636 2465
rect 25044 2456 25096 2508
rect 25228 2499 25280 2508
rect 25228 2465 25237 2499
rect 25237 2465 25271 2499
rect 25271 2465 25280 2499
rect 25228 2456 25280 2465
rect 6460 2320 6512 2372
rect 8852 2320 8904 2372
rect 13820 2388 13872 2440
rect 14096 2388 14148 2440
rect 15384 2320 15436 2372
rect 16856 2320 16908 2372
rect 18788 2320 18840 2372
rect 21364 2320 21416 2372
rect 14280 2252 14332 2304
rect 28816 2524 28868 2576
rect 29736 2524 29788 2576
rect 27620 2456 27672 2508
rect 27804 2499 27856 2508
rect 27804 2465 27813 2499
rect 27813 2465 27847 2499
rect 27847 2465 27856 2499
rect 27804 2456 27856 2465
rect 30748 2456 30800 2508
rect 32220 2524 32272 2576
rect 31944 2456 31996 2508
rect 37556 2524 37608 2576
rect 32404 2456 32456 2508
rect 34244 2456 34296 2508
rect 37280 2499 37332 2508
rect 37280 2465 37289 2499
rect 37289 2465 37323 2499
rect 37323 2465 37332 2499
rect 37280 2456 37332 2465
rect 38292 2456 38344 2508
rect 39488 2524 39540 2576
rect 39396 2456 39448 2508
rect 40040 2499 40092 2508
rect 40040 2465 40049 2499
rect 40049 2465 40083 2499
rect 40083 2465 40092 2499
rect 40040 2456 40092 2465
rect 43536 2524 43588 2576
rect 44548 2524 44600 2576
rect 42616 2499 42668 2508
rect 42616 2465 42625 2499
rect 42625 2465 42659 2499
rect 42659 2465 42668 2499
rect 42616 2456 42668 2465
rect 42708 2456 42760 2508
rect 45560 2456 45612 2508
rect 34704 2431 34756 2440
rect 34704 2397 34713 2431
rect 34713 2397 34747 2431
rect 34747 2397 34756 2431
rect 34704 2388 34756 2397
rect 29092 2320 29144 2372
rect 34520 2320 34572 2372
rect 44456 2320 44508 2372
rect 38476 2252 38528 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 14004 1504 14056 1556
rect 14924 1504 14976 1556
<< metal2 >>
rect 1738 49200 1850 50000
rect 5050 49314 5162 50000
rect 5050 49286 5304 49314
rect 5050 49200 5162 49286
rect 1780 47054 1808 49200
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 2228 47184 2280 47190
rect 2228 47126 2280 47132
rect 1768 47048 1820 47054
rect 1768 46990 1820 46996
rect 2240 16574 2268 47126
rect 5276 47054 5304 49286
rect 8362 49200 8474 50000
rect 11674 49200 11786 50000
rect 14986 49200 15098 50000
rect 18298 49200 18410 50000
rect 21610 49314 21722 50000
rect 21610 49286 21864 49314
rect 21610 49200 21722 49286
rect 21836 47054 21864 49286
rect 24922 49200 25034 50000
rect 28234 49200 28346 50000
rect 31546 49200 31658 50000
rect 34858 49200 34970 50000
rect 38170 49200 38282 50000
rect 41482 49200 41594 50000
rect 44794 49200 44906 50000
rect 48106 49200 48218 50000
rect 24964 47054 24992 49200
rect 28276 47054 28304 49200
rect 31588 47138 31616 49200
rect 34900 47546 34928 49200
rect 34808 47518 34928 47546
rect 31588 47110 31800 47138
rect 31772 47054 31800 47110
rect 34808 47054 34836 47518
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34888 47184 34940 47190
rect 34888 47126 34940 47132
rect 5264 47048 5316 47054
rect 5264 46990 5316 46996
rect 21824 47048 21876 47054
rect 21824 46990 21876 46996
rect 24952 47048 25004 47054
rect 24952 46990 25004 46996
rect 28264 47048 28316 47054
rect 28264 46990 28316 46996
rect 31760 47048 31812 47054
rect 31760 46990 31812 46996
rect 34796 47048 34848 47054
rect 34796 46990 34848 46996
rect 8208 46980 8260 46986
rect 8208 46922 8260 46928
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 2240 16546 2360 16574
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 756 4004 808 4010
rect 756 3946 808 3952
rect 768 800 796 3946
rect 1412 2514 1440 7890
rect 1596 4146 1624 8298
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1596 1714 1624 3538
rect 1688 2514 1716 6054
rect 1780 4078 1808 7142
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1872 3738 1900 7822
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1964 6798 1992 7346
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1964 6322 1992 6734
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 2056 3466 2084 6598
rect 2332 5234 2360 16546
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2608 5302 2636 6258
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 2240 4282 2268 4422
rect 2228 4276 2280 4282
rect 2228 4218 2280 4224
rect 2332 4214 2360 5170
rect 2700 4622 2728 5170
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2320 4208 2372 4214
rect 2320 4150 2372 4156
rect 2044 3460 2096 3466
rect 2044 3402 2096 3408
rect 2792 3194 2820 7142
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2884 4690 2912 5102
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2872 4548 2924 4554
rect 2872 4490 2924 4496
rect 2884 3670 2912 4490
rect 3068 4185 3096 4966
rect 3054 4176 3110 4185
rect 3054 4111 3110 4120
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 3160 3126 3188 6598
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3252 4690 3280 5714
rect 3344 5710 3372 6734
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 3698 6352 3754 6361
rect 3698 6287 3754 6296
rect 4068 6316 4120 6322
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3148 3120 3200 3126
rect 3148 3062 3200 3068
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 1412 1686 1624 1714
rect 1412 800 1440 1686
rect 2056 800 2084 2450
rect 2700 800 2728 2926
rect 3344 800 3372 3946
rect 3436 2514 3464 6054
rect 3620 4554 3648 6122
rect 3712 5710 3740 6287
rect 4068 6258 4120 6264
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3700 5704 3752 5710
rect 3988 5681 4016 6054
rect 3700 5646 3752 5652
rect 3974 5672 4030 5681
rect 3712 5234 3740 5646
rect 3974 5607 4030 5616
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3608 4548 3660 4554
rect 3608 4490 3660 4496
rect 3804 4078 3832 5510
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3988 4146 4016 5034
rect 4080 4826 4108 6258
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5896 4660 6666
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4540 5868 4660 5896
rect 4436 5704 4488 5710
rect 4540 5692 4568 5868
rect 4488 5664 4568 5692
rect 4618 5672 4674 5681
rect 4436 5646 4488 5652
rect 4252 5636 4304 5642
rect 4618 5607 4620 5616
rect 4252 5578 4304 5584
rect 4672 5607 4674 5616
rect 4620 5578 4672 5584
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4172 5370 4200 5510
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4264 5114 4292 5578
rect 4264 5086 4660 5114
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 4264 4010 4292 4626
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3988 800 4016 3878
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3126 4660 5086
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4724 2774 4752 6598
rect 4816 2990 4844 6734
rect 5000 6662 5028 7346
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 5092 7002 5120 7142
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5000 6322 5028 6598
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 4988 6180 5040 6186
rect 4988 6122 5040 6128
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4908 4758 4936 6054
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 5000 3670 5028 6122
rect 5092 5302 5120 6394
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 4988 3664 5040 3670
rect 4988 3606 5040 3612
rect 5184 3602 5212 7686
rect 6104 7410 6132 7822
rect 7668 7818 7696 8434
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6644 7404 6696 7410
rect 6696 7364 6776 7392
rect 6644 7346 6696 7352
rect 5552 6866 5580 7346
rect 6368 7268 6420 7274
rect 6368 7210 6420 7216
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5264 6316 5316 6322
rect 5316 6276 5580 6304
rect 5264 6258 5316 6264
rect 5552 5166 5580 6276
rect 5644 5234 5672 6598
rect 5736 6322 5764 6666
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5552 4690 5580 5102
rect 5828 5098 5856 6802
rect 6380 6322 6408 7210
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 6196 4690 6224 5510
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 5552 4282 5580 4626
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 5264 2916 5316 2922
rect 5264 2858 5316 2864
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2746 4752 2774
rect 4632 2650 4660 2746
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4632 800 4660 2450
rect 5276 800 5304 2858
rect 5920 800 5948 3538
rect 6288 3466 6316 5850
rect 6380 5710 6408 6258
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6472 4690 6500 7142
rect 6748 6254 6776 7364
rect 7116 6730 7144 7686
rect 7208 7410 7236 7754
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6656 5370 6684 6190
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6840 5370 6868 5510
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 7116 5302 7144 6054
rect 7300 5778 7328 7142
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7576 5778 7604 6666
rect 7760 6322 7788 8298
rect 8220 7886 8248 46922
rect 22008 46912 22060 46918
rect 22008 46854 22060 46860
rect 25228 46912 25280 46918
rect 25228 46854 25280 46860
rect 28540 46912 28592 46918
rect 28540 46854 28592 46860
rect 32312 46912 32364 46918
rect 32312 46854 32364 46860
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8496 7478 8524 8026
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8036 6458 8064 6598
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8128 6361 8156 6394
rect 8114 6352 8170 6361
rect 7748 6316 7800 6322
rect 8114 6287 8170 6296
rect 7748 6258 7800 6264
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7208 5370 7236 5510
rect 7576 5370 7604 5714
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7104 5296 7156 5302
rect 7104 5238 7156 5244
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6276 3460 6328 3466
rect 6276 3402 6328 3408
rect 6472 2378 6500 4422
rect 6564 2514 6592 5102
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6932 2774 6960 4626
rect 7010 4176 7066 4185
rect 7010 4111 7066 4120
rect 7024 4078 7052 4111
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 7116 4010 7144 5238
rect 7208 5166 7236 5306
rect 8404 5302 8432 5782
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8496 5166 8524 7414
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8680 5710 8708 6054
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 6656 2746 6960 2774
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 6460 2372 6512 2378
rect 6460 2314 6512 2320
rect 6656 1442 6684 2746
rect 6564 1414 6684 1442
rect 6564 800 6592 1414
rect 7208 800 7236 4014
rect 8484 3460 8536 3466
rect 8484 3402 8536 3408
rect 7748 2508 7800 2514
rect 7800 2468 7880 2496
rect 7748 2450 7800 2456
rect 7852 800 7880 2468
rect 8496 800 8524 3402
rect 8864 2378 8892 8298
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 8956 6798 8984 7754
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8956 6322 8984 6734
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 9048 3126 9076 8298
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9140 5302 9168 6598
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9232 4690 9260 7686
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9324 4078 9352 8298
rect 9600 7886 9628 8366
rect 10336 7954 10364 8910
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9508 6866 9536 7278
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9416 6186 9444 6734
rect 9600 6458 9628 7822
rect 10232 7812 10284 7818
rect 10232 7754 10284 7760
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9508 5710 9536 6258
rect 9692 5778 9720 6258
rect 9784 6254 9812 6734
rect 9876 6390 9904 7142
rect 10244 6866 10272 7754
rect 10428 7478 10456 8774
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10980 7886 11008 8434
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10416 7472 10468 7478
rect 10416 7414 10468 7420
rect 10980 7410 11008 7822
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 10244 5914 10272 6326
rect 10336 6322 10364 6598
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9508 5030 9536 5646
rect 9600 5302 9628 5646
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9508 3670 9536 4966
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 9600 3602 9628 5238
rect 10244 5234 10272 5850
rect 10336 5370 10364 6258
rect 10612 6254 10640 6666
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10520 5574 10548 5714
rect 10508 5568 10560 5574
rect 10508 5510 10560 5516
rect 10520 5370 10548 5510
rect 10704 5370 10732 5714
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 9140 800 9168 2450
rect 9784 800 9812 4626
rect 10244 2582 10272 5170
rect 10336 4758 10364 5306
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10232 2576 10284 2582
rect 10232 2518 10284 2524
rect 10428 800 10456 3538
rect 11072 2990 11100 7686
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11164 3466 11192 7210
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11440 3466 11468 7142
rect 11900 6730 11928 8774
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 12452 6458 12480 7346
rect 12544 6798 12572 8910
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 22020 6914 22048 46854
rect 21744 6886 22048 6914
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11808 5914 11836 6122
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 12360 5846 12388 6258
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12452 5914 12480 6054
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12348 5840 12400 5846
rect 12348 5782 12400 5788
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 11808 5302 11836 5714
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 11072 800 11100 2790
rect 11716 800 11744 4014
rect 12176 2990 12204 5578
rect 12452 4554 12480 5714
rect 13188 5302 13216 6598
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 13452 6180 13504 6186
rect 13452 6122 13504 6128
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 13464 4078 13492 6122
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13636 4548 13688 4554
rect 13636 4490 13688 4496
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13096 3942 13124 4014
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 13280 3738 13308 4014
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 12992 3460 13044 3466
rect 12992 3402 13044 3408
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 12164 2984 12216 2990
rect 11900 2922 12112 2938
rect 12164 2926 12216 2932
rect 11888 2916 12124 2922
rect 11940 2910 12072 2916
rect 11888 2858 11940 2864
rect 12072 2858 12124 2864
rect 12360 800 12388 3062
rect 13004 800 13032 3402
rect 13648 800 13676 4490
rect 13832 2446 13860 6054
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 13924 4214 13952 5782
rect 14384 5710 14412 6258
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14096 5092 14148 5098
rect 14096 5034 14148 5040
rect 13912 4208 13964 4214
rect 13912 4150 13964 4156
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 14016 1562 14044 2926
rect 14108 2446 14136 5034
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14384 3602 14412 4966
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14476 3466 14504 5510
rect 14936 4758 14964 5646
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 21088 5228 21140 5234
rect 21088 5170 21140 5176
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 14648 4548 14700 4554
rect 14648 4490 14700 4496
rect 14660 4214 14688 4490
rect 14648 4208 14700 4214
rect 14648 4150 14700 4156
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14200 3058 14228 3334
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 15212 2990 15240 4966
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15200 2984 15252 2990
rect 14200 2922 14596 2938
rect 15200 2926 15252 2932
rect 14188 2916 14608 2922
rect 14240 2910 14556 2916
rect 14188 2858 14240 2864
rect 14556 2858 14608 2864
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 15396 2378 15424 4422
rect 15856 4146 15884 4558
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14004 1556 14056 1562
rect 14004 1498 14056 1504
rect 14292 800 14320 2246
rect 14924 1556 14976 1562
rect 14924 1498 14976 1504
rect 14936 800 14964 1498
rect 15580 800 15608 4014
rect 15948 3398 15976 4966
rect 16120 4616 16172 4622
rect 16120 4558 16172 4564
rect 16132 3602 16160 4558
rect 16500 4146 16528 5170
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 16316 3466 16344 3878
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 16224 800 16252 3402
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16684 3194 16712 3334
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16776 2514 16804 4558
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 17052 2514 17080 3878
rect 17144 3058 17172 4558
rect 17420 3602 17448 4966
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 17500 3120 17552 3126
rect 17500 3062 17552 3068
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 16764 2508 16816 2514
rect 16764 2450 16816 2456
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 16856 2372 16908 2378
rect 16856 2314 16908 2320
rect 16868 800 16896 2314
rect 17512 800 17540 3062
rect 17972 2990 18000 4966
rect 18432 4622 18460 5170
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18064 4146 18092 4558
rect 18432 4214 18460 4558
rect 18696 4480 18748 4486
rect 18696 4422 18748 4428
rect 18708 4214 18736 4422
rect 18420 4208 18472 4214
rect 18420 4150 18472 4156
rect 18696 4208 18748 4214
rect 18696 4150 18748 4156
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 19168 3602 19196 4966
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 18156 800 18184 3538
rect 19352 2514 19380 4966
rect 19432 4548 19484 4554
rect 19432 4490 19484 4496
rect 19444 4162 19472 4490
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19444 4134 19564 4162
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19444 3602 19472 3878
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19536 3466 19564 4134
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 18788 2372 18840 2378
rect 18788 2314 18840 2320
rect 18800 800 18828 2314
rect 19444 800 19472 3062
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 20088 800 20116 4014
rect 20364 2514 20392 4966
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20548 4282 20576 4558
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 20732 800 20760 3538
rect 20824 2990 20852 4966
rect 21100 4554 21128 5170
rect 21456 5024 21508 5030
rect 21456 4966 21508 4972
rect 21088 4548 21140 4554
rect 21088 4490 21140 4496
rect 21100 4214 21128 4490
rect 21088 4208 21140 4214
rect 21088 4150 21140 4156
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 21376 2854 21404 3130
rect 21468 3126 21496 4966
rect 21744 3398 21772 6886
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 23848 5024 23900 5030
rect 23848 4966 23900 4972
rect 24584 5024 24636 5030
rect 24584 4966 24636 4972
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 21928 3602 21956 4558
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21732 3392 21784 3398
rect 21732 3334 21784 3340
rect 21456 3120 21508 3126
rect 21456 3062 21508 3068
rect 21916 2984 21968 2990
rect 21916 2926 21968 2932
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21364 2372 21416 2378
rect 21364 2314 21416 2320
rect 21376 800 21404 2314
rect 21928 1578 21956 2926
rect 22020 2514 22048 3878
rect 22112 3466 22140 4422
rect 22100 3460 22152 3466
rect 22100 3402 22152 3408
rect 22296 3058 22324 4966
rect 23296 4616 23348 4622
rect 23296 4558 23348 4564
rect 23112 4480 23164 4486
rect 23112 4422 23164 4428
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22480 3126 22508 3878
rect 22652 3460 22704 3466
rect 22652 3402 22704 3408
rect 22468 3120 22520 3126
rect 22468 3062 22520 3068
rect 22284 3052 22336 3058
rect 22284 2994 22336 3000
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 21928 1550 22048 1578
rect 22020 800 22048 1550
rect 22664 800 22692 3402
rect 23124 2514 23152 4422
rect 23308 4282 23336 4558
rect 23388 4548 23440 4554
rect 23388 4490 23440 4496
rect 23296 4276 23348 4282
rect 23296 4218 23348 4224
rect 23308 4078 23336 4218
rect 23400 4214 23428 4490
rect 23388 4208 23440 4214
rect 23388 4150 23440 4156
rect 23860 4146 23888 4966
rect 24032 4480 24084 4486
rect 24032 4422 24084 4428
rect 24044 4214 24072 4422
rect 24032 4208 24084 4214
rect 24032 4150 24084 4156
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 24492 4072 24544 4078
rect 24492 4014 24544 4020
rect 23940 2984 23992 2990
rect 23940 2926 23992 2932
rect 23112 2508 23164 2514
rect 23112 2450 23164 2456
rect 23388 2508 23440 2514
rect 23388 2450 23440 2456
rect 23400 1170 23428 2450
rect 23308 1142 23428 1170
rect 23308 800 23336 1142
rect 23952 800 23980 2926
rect 24504 2122 24532 4014
rect 24596 2514 24624 4966
rect 24952 4752 25004 4758
rect 24952 4694 25004 4700
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24780 3126 24808 4422
rect 24964 3670 24992 4694
rect 25240 4010 25268 46854
rect 28552 6914 28580 46854
rect 32324 16574 32352 46854
rect 34900 46458 34928 47126
rect 38212 47054 38240 49200
rect 38200 47048 38252 47054
rect 38200 46990 38252 46996
rect 41524 46918 41552 49200
rect 44836 47054 44864 49200
rect 48148 47054 48176 49200
rect 44824 47048 44876 47054
rect 44824 46990 44876 46996
rect 48136 47048 48188 47054
rect 48136 46990 48188 46996
rect 47952 46980 48004 46986
rect 47952 46922 48004 46928
rect 38476 46912 38528 46918
rect 38476 46854 38528 46860
rect 41512 46912 41564 46918
rect 41512 46854 41564 46860
rect 42984 46912 43036 46918
rect 42984 46854 43036 46860
rect 45560 46912 45612 46918
rect 45560 46854 45612 46860
rect 34808 46430 34928 46458
rect 32324 16546 32536 16574
rect 28368 6886 28580 6914
rect 25320 4616 25372 4622
rect 25320 4558 25372 4564
rect 27620 4616 27672 4622
rect 27620 4558 27672 4564
rect 25228 4004 25280 4010
rect 25228 3946 25280 3952
rect 24952 3664 25004 3670
rect 24952 3606 25004 3612
rect 24964 3534 24992 3606
rect 24952 3528 25004 3534
rect 24952 3470 25004 3476
rect 25044 3392 25096 3398
rect 25044 3334 25096 3340
rect 24768 3120 24820 3126
rect 24768 3062 24820 3068
rect 25056 2514 25084 3334
rect 25332 2990 25360 4558
rect 25872 4480 25924 4486
rect 25872 4422 25924 4428
rect 25688 3936 25740 3942
rect 25688 3878 25740 3884
rect 25700 3534 25728 3878
rect 25688 3528 25740 3534
rect 25688 3470 25740 3476
rect 25884 3466 25912 4422
rect 27632 4146 27660 4558
rect 27620 4140 27672 4146
rect 27620 4082 27672 4088
rect 27632 4026 27660 4082
rect 26240 4004 26292 4010
rect 27632 3998 27752 4026
rect 26240 3946 26292 3952
rect 26252 3602 26280 3946
rect 26976 3936 27028 3942
rect 26976 3878 27028 3884
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 26240 3596 26292 3602
rect 26240 3538 26292 3544
rect 26516 3596 26568 3602
rect 26516 3538 26568 3544
rect 25872 3460 25924 3466
rect 25872 3402 25924 3408
rect 25320 2984 25372 2990
rect 25320 2926 25372 2932
rect 25964 2984 26016 2990
rect 25964 2926 26016 2932
rect 24584 2508 24636 2514
rect 24584 2450 24636 2456
rect 25044 2508 25096 2514
rect 25044 2450 25096 2456
rect 25228 2508 25280 2514
rect 25228 2450 25280 2456
rect 24504 2094 24624 2122
rect 24596 800 24624 2094
rect 25240 800 25268 2450
rect 25976 1578 26004 2926
rect 25884 1550 26004 1578
rect 25884 800 25912 1550
rect 26528 800 26556 3538
rect 26988 3058 27016 3878
rect 27160 3392 27212 3398
rect 27160 3334 27212 3340
rect 27172 3126 27200 3334
rect 27160 3120 27212 3126
rect 27160 3062 27212 3068
rect 26976 3052 27028 3058
rect 26976 2994 27028 3000
rect 27160 2984 27212 2990
rect 27160 2926 27212 2932
rect 27172 800 27200 2926
rect 27632 2514 27660 3878
rect 27724 3534 27752 3998
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 28368 2854 28396 6886
rect 31852 5772 31904 5778
rect 31852 5714 31904 5720
rect 28540 5228 28592 5234
rect 28540 5170 28592 5176
rect 31668 5228 31720 5234
rect 31668 5170 31720 5176
rect 28448 5024 28500 5030
rect 28448 4966 28500 4972
rect 28460 4214 28488 4966
rect 28552 4622 28580 5170
rect 29092 5024 29144 5030
rect 29092 4966 29144 4972
rect 28908 4684 28960 4690
rect 28908 4626 28960 4632
rect 28540 4616 28592 4622
rect 28540 4558 28592 4564
rect 28448 4208 28500 4214
rect 28448 4150 28500 4156
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 28448 2848 28500 2854
rect 28448 2790 28500 2796
rect 27620 2508 27672 2514
rect 27620 2450 27672 2456
rect 27804 2508 27856 2514
rect 27804 2450 27856 2456
rect 27816 800 27844 2450
rect 28460 800 28488 2790
rect 28828 2582 28856 3470
rect 28920 3058 28948 4626
rect 28908 3052 28960 3058
rect 28908 2994 28960 3000
rect 28816 2576 28868 2582
rect 28816 2518 28868 2524
rect 29104 2378 29132 4966
rect 31680 4826 31708 5170
rect 31668 4820 31720 4826
rect 31668 4762 31720 4768
rect 29736 4616 29788 4622
rect 29736 4558 29788 4564
rect 30380 4616 30432 4622
rect 30380 4558 30432 4564
rect 29460 4480 29512 4486
rect 29460 4422 29512 4428
rect 29184 4004 29236 4010
rect 29184 3946 29236 3952
rect 29092 2372 29144 2378
rect 29092 2314 29144 2320
rect 29196 2122 29224 3946
rect 29472 3126 29500 4422
rect 29748 4078 29776 4558
rect 29736 4072 29788 4078
rect 29736 4014 29788 4020
rect 30392 3670 30420 4558
rect 31680 4146 31708 4762
rect 31760 4616 31812 4622
rect 31760 4558 31812 4564
rect 31668 4140 31720 4146
rect 31668 4082 31720 4088
rect 30748 3936 30800 3942
rect 30748 3878 30800 3884
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 30380 3664 30432 3670
rect 30380 3606 30432 3612
rect 30380 3460 30432 3466
rect 30380 3402 30432 3408
rect 29460 3120 29512 3126
rect 29460 3062 29512 3068
rect 29736 2576 29788 2582
rect 29736 2518 29788 2524
rect 29104 2094 29224 2122
rect 29104 800 29132 2094
rect 29748 800 29776 2518
rect 30392 800 30420 3402
rect 30760 2514 30788 3878
rect 31312 3602 31340 3878
rect 31668 3664 31720 3670
rect 31668 3606 31720 3612
rect 31300 3596 31352 3602
rect 31300 3538 31352 3544
rect 31024 2848 31076 2854
rect 31024 2790 31076 2796
rect 30748 2508 30800 2514
rect 30748 2450 30800 2456
rect 31036 800 31064 2790
rect 31680 800 31708 3606
rect 31772 3058 31800 4558
rect 31864 3602 31892 5714
rect 31944 5704 31996 5710
rect 31944 5646 31996 5652
rect 32128 5704 32180 5710
rect 32128 5646 32180 5652
rect 31852 3596 31904 3602
rect 31852 3538 31904 3544
rect 31760 3052 31812 3058
rect 31760 2994 31812 3000
rect 31956 2514 31984 5646
rect 32036 5024 32088 5030
rect 32036 4966 32088 4972
rect 32048 3602 32076 4966
rect 32140 4146 32168 5646
rect 32404 5092 32456 5098
rect 32404 5034 32456 5040
rect 32220 5024 32272 5030
rect 32220 4966 32272 4972
rect 32312 5024 32364 5030
rect 32312 4966 32364 4972
rect 32128 4140 32180 4146
rect 32128 4082 32180 4088
rect 32036 3596 32088 3602
rect 32036 3538 32088 3544
rect 32232 2582 32260 4966
rect 32324 4214 32352 4966
rect 32312 4208 32364 4214
rect 32312 4150 32364 4156
rect 32416 3126 32444 5034
rect 32508 4010 32536 16546
rect 33416 5228 33468 5234
rect 33416 5170 33468 5176
rect 33428 4826 33456 5170
rect 34612 5092 34664 5098
rect 34612 5034 34664 5040
rect 34520 5024 34572 5030
rect 34520 4966 34572 4972
rect 33416 4820 33468 4826
rect 33416 4762 33468 4768
rect 34428 4616 34480 4622
rect 34428 4558 34480 4564
rect 32956 4072 33008 4078
rect 32956 4014 33008 4020
rect 32496 4004 32548 4010
rect 32496 3946 32548 3952
rect 32404 3120 32456 3126
rect 32404 3062 32456 3068
rect 32220 2576 32272 2582
rect 32220 2518 32272 2524
rect 31944 2508 31996 2514
rect 31944 2450 31996 2456
rect 32404 2508 32456 2514
rect 32404 2450 32456 2456
rect 32416 1170 32444 2450
rect 32324 1142 32444 1170
rect 32324 800 32352 1142
rect 32968 800 32996 4014
rect 34440 3058 34468 4558
rect 33600 3052 33652 3058
rect 33600 2994 33652 3000
rect 34428 3052 34480 3058
rect 34428 2994 34480 3000
rect 33612 800 33640 2994
rect 34244 2508 34296 2514
rect 34244 2450 34296 2456
rect 34256 800 34284 2450
rect 34532 2378 34560 4966
rect 34624 3126 34652 5034
rect 34704 5024 34756 5030
rect 34704 4966 34756 4972
rect 34716 3602 34744 4966
rect 34808 4758 34836 46430
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 36360 5704 36412 5710
rect 36360 5646 36412 5652
rect 37280 5704 37332 5710
rect 37280 5646 37332 5652
rect 35440 5228 35492 5234
rect 35440 5170 35492 5176
rect 35348 5024 35400 5030
rect 35348 4966 35400 4972
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34796 4752 34848 4758
rect 34796 4694 34848 4700
rect 34796 4616 34848 4622
rect 34796 4558 34848 4564
rect 34704 3596 34756 3602
rect 34704 3538 34756 3544
rect 34808 3482 34836 4558
rect 35360 4214 35388 4966
rect 35452 4622 35480 5170
rect 35440 4616 35492 4622
rect 35440 4558 35492 4564
rect 36176 4616 36228 4622
rect 36176 4558 36228 4564
rect 35440 4480 35492 4486
rect 35440 4422 35492 4428
rect 35348 4208 35400 4214
rect 35348 4150 35400 4156
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34888 3596 34940 3602
rect 34888 3538 34940 3544
rect 34716 3454 34836 3482
rect 34612 3120 34664 3126
rect 34612 3062 34664 3068
rect 34716 2446 34744 3454
rect 34900 2904 34928 3538
rect 35452 3466 35480 4422
rect 36188 4078 36216 4558
rect 36176 4072 36228 4078
rect 36176 4014 36228 4020
rect 35532 4004 35584 4010
rect 35532 3946 35584 3952
rect 35440 3460 35492 3466
rect 35440 3402 35492 3408
rect 34808 2876 34928 2904
rect 34704 2440 34756 2446
rect 34704 2382 34756 2388
rect 34520 2372 34572 2378
rect 34520 2314 34572 2320
rect 34808 1850 34836 2876
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34808 1822 34928 1850
rect 34900 800 34928 1822
rect 35544 800 35572 3946
rect 36372 3602 36400 5646
rect 36820 3664 36872 3670
rect 36820 3606 36872 3612
rect 36360 3596 36412 3602
rect 36360 3538 36412 3544
rect 36176 2916 36228 2922
rect 36176 2858 36228 2864
rect 36188 800 36216 2858
rect 36832 800 36860 3606
rect 37292 2514 37320 5646
rect 37924 5228 37976 5234
rect 37924 5170 37976 5176
rect 37648 5092 37700 5098
rect 37648 5034 37700 5040
rect 37372 5024 37424 5030
rect 37372 4966 37424 4972
rect 37556 5024 37608 5030
rect 37556 4966 37608 4972
rect 37384 3602 37412 4966
rect 37464 4480 37516 4486
rect 37464 4422 37516 4428
rect 37372 3596 37424 3602
rect 37372 3538 37424 3544
rect 37476 3126 37504 4422
rect 37568 4214 37596 4966
rect 37556 4208 37608 4214
rect 37556 4150 37608 4156
rect 37464 3120 37516 3126
rect 37464 3062 37516 3068
rect 37660 2990 37688 5034
rect 37936 4622 37964 5170
rect 37924 4616 37976 4622
rect 37924 4558 37976 4564
rect 37740 4480 37792 4486
rect 37740 4422 37792 4428
rect 38292 4480 38344 4486
rect 38292 4422 38344 4428
rect 37752 3398 37780 4422
rect 38108 4072 38160 4078
rect 38108 4014 38160 4020
rect 37740 3392 37792 3398
rect 37740 3334 37792 3340
rect 37648 2984 37700 2990
rect 37648 2926 37700 2932
rect 37556 2576 37608 2582
rect 37556 2518 37608 2524
rect 37280 2508 37332 2514
rect 37280 2450 37332 2456
rect 37568 1170 37596 2518
rect 37476 1142 37596 1170
rect 37476 800 37504 1142
rect 38120 800 38148 4014
rect 38304 2514 38332 4422
rect 38292 2508 38344 2514
rect 38292 2450 38344 2456
rect 38488 2310 38516 46854
rect 39580 5704 39632 5710
rect 39580 5646 39632 5652
rect 40132 5704 40184 5710
rect 40132 5646 40184 5652
rect 41604 5704 41656 5710
rect 41604 5646 41656 5652
rect 38660 5024 38712 5030
rect 38660 4966 38712 4972
rect 39396 5024 39448 5030
rect 39396 4966 39448 4972
rect 38672 3126 38700 4966
rect 39028 4616 39080 4622
rect 39028 4558 39080 4564
rect 39040 4010 39068 4558
rect 39028 4004 39080 4010
rect 39028 3946 39080 3952
rect 38660 3120 38712 3126
rect 38660 3062 38712 3068
rect 38752 2984 38804 2990
rect 38752 2926 38804 2932
rect 38476 2304 38528 2310
rect 38476 2246 38528 2252
rect 38764 800 38792 2926
rect 39408 2514 39436 4966
rect 39592 3058 39620 5646
rect 40040 4480 40092 4486
rect 40040 4422 40092 4428
rect 39580 3052 39632 3058
rect 39580 2994 39632 3000
rect 39488 2576 39540 2582
rect 39488 2518 39540 2524
rect 39396 2508 39448 2514
rect 39396 2450 39448 2456
rect 39500 1170 39528 2518
rect 40052 2514 40080 4422
rect 40144 4010 40172 5646
rect 40224 5024 40276 5030
rect 40224 4966 40276 4972
rect 40592 5024 40644 5030
rect 40592 4966 40644 4972
rect 40132 4004 40184 4010
rect 40132 3946 40184 3952
rect 40132 3664 40184 3670
rect 40132 3606 40184 3612
rect 40040 2508 40092 2514
rect 40040 2450 40092 2456
rect 40144 1714 40172 3606
rect 40236 3602 40264 4966
rect 40224 3596 40276 3602
rect 40224 3538 40276 3544
rect 40604 3466 40632 4966
rect 41512 4480 41564 4486
rect 41512 4422 41564 4428
rect 41524 4078 41552 4422
rect 41512 4072 41564 4078
rect 41512 4014 41564 4020
rect 40684 4004 40736 4010
rect 40684 3946 40736 3952
rect 40592 3460 40644 3466
rect 40592 3402 40644 3408
rect 39408 1142 39528 1170
rect 40052 1686 40172 1714
rect 39408 800 39436 1142
rect 40052 800 40080 1686
rect 40696 800 40724 3946
rect 41616 3602 41644 5646
rect 42432 5228 42484 5234
rect 42432 5170 42484 5176
rect 42064 5024 42116 5030
rect 42064 4966 42116 4972
rect 41972 3664 42024 3670
rect 41972 3606 42024 3612
rect 41604 3596 41656 3602
rect 41604 3538 41656 3544
rect 41328 2984 41380 2990
rect 41328 2926 41380 2932
rect 41340 800 41368 2926
rect 41984 800 42012 3606
rect 42076 3126 42104 4966
rect 42444 4622 42472 5170
rect 42616 5024 42668 5030
rect 42616 4966 42668 4972
rect 42248 4616 42300 4622
rect 42248 4558 42300 4564
rect 42432 4616 42484 4622
rect 42432 4558 42484 4564
rect 42064 3120 42116 3126
rect 42064 3062 42116 3068
rect 42260 3058 42288 4558
rect 42248 3052 42300 3058
rect 42248 2994 42300 3000
rect 42628 2514 42656 4966
rect 42800 4480 42852 4486
rect 42800 4422 42852 4428
rect 42812 3602 42840 4422
rect 42800 3596 42852 3602
rect 42800 3538 42852 3544
rect 42996 2854 43024 46854
rect 45376 8356 45428 8362
rect 45376 8298 45428 8304
rect 45284 7336 45336 7342
rect 45284 7278 45336 7284
rect 45008 5704 45060 5710
rect 45008 5646 45060 5652
rect 44916 5568 44968 5574
rect 44916 5510 44968 5516
rect 43260 5024 43312 5030
rect 43260 4966 43312 4972
rect 43812 5024 43864 5030
rect 43812 4966 43864 4972
rect 44456 5024 44508 5030
rect 44456 4966 44508 4972
rect 43272 4214 43300 4966
rect 43536 4616 43588 4622
rect 43536 4558 43588 4564
rect 43260 4208 43312 4214
rect 43260 4150 43312 4156
rect 43260 4004 43312 4010
rect 43260 3946 43312 3952
rect 42984 2848 43036 2854
rect 42984 2790 43036 2796
rect 42616 2508 42668 2514
rect 42616 2450 42668 2456
rect 42708 2508 42760 2514
rect 42708 2450 42760 2456
rect 42720 1170 42748 2450
rect 42628 1142 42748 1170
rect 42628 800 42656 1142
rect 43272 800 43300 3946
rect 43548 2582 43576 4558
rect 43824 4078 43852 4966
rect 43812 4072 43864 4078
rect 43812 4014 43864 4020
rect 43904 2848 43956 2854
rect 43904 2790 43956 2796
rect 43536 2576 43588 2582
rect 43536 2518 43588 2524
rect 43916 800 43944 2790
rect 44468 2378 44496 4966
rect 44928 3126 44956 5510
rect 45020 5234 45048 5646
rect 45192 5568 45244 5574
rect 45192 5510 45244 5516
rect 45008 5228 45060 5234
rect 45008 5170 45060 5176
rect 45020 4554 45048 5170
rect 45008 4548 45060 4554
rect 45008 4490 45060 4496
rect 45204 4078 45232 5510
rect 45296 5250 45324 7278
rect 45388 6254 45416 8298
rect 45468 7268 45520 7274
rect 45468 7210 45520 7216
rect 45376 6248 45428 6254
rect 45376 6190 45428 6196
rect 45480 5302 45508 7210
rect 45468 5296 45520 5302
rect 45296 5222 45416 5250
rect 45468 5238 45520 5244
rect 45388 5166 45416 5222
rect 45376 5160 45428 5166
rect 45376 5102 45428 5108
rect 45376 4548 45428 4554
rect 45376 4490 45428 4496
rect 45192 4072 45244 4078
rect 45192 4014 45244 4020
rect 45388 3738 45416 4490
rect 45376 3732 45428 3738
rect 45376 3674 45428 3680
rect 45572 3670 45600 46854
rect 47584 8492 47636 8498
rect 47584 8434 47636 8440
rect 47596 7886 47624 8434
rect 47124 7880 47176 7886
rect 47124 7822 47176 7828
rect 47584 7880 47636 7886
rect 47584 7822 47636 7828
rect 46388 7200 46440 7206
rect 46388 7142 46440 7148
rect 46400 6390 46428 7142
rect 47136 6866 47164 7822
rect 47596 7410 47624 7822
rect 47964 7818 47992 46922
rect 47952 7812 48004 7818
rect 47952 7754 48004 7760
rect 47676 7744 47728 7750
rect 47676 7686 47728 7692
rect 47584 7404 47636 7410
rect 47584 7346 47636 7352
rect 47124 6860 47176 6866
rect 47124 6802 47176 6808
rect 46388 6384 46440 6390
rect 46388 6326 46440 6332
rect 46296 6112 46348 6118
rect 46296 6054 46348 6060
rect 46308 5778 46336 6054
rect 45836 5772 45888 5778
rect 45836 5714 45888 5720
rect 46296 5772 46348 5778
rect 46296 5714 46348 5720
rect 47124 5772 47176 5778
rect 47124 5714 47176 5720
rect 45652 5704 45704 5710
rect 45652 5646 45704 5652
rect 45664 5166 45692 5646
rect 45652 5160 45704 5166
rect 45652 5102 45704 5108
rect 45664 4826 45692 5102
rect 45652 4820 45704 4826
rect 45652 4762 45704 4768
rect 45848 4690 45876 5714
rect 46020 5024 46072 5030
rect 46020 4966 46072 4972
rect 46032 4690 46060 4966
rect 45836 4684 45888 4690
rect 45836 4626 45888 4632
rect 46020 4684 46072 4690
rect 46020 4626 46072 4632
rect 46480 4684 46532 4690
rect 46480 4626 46532 4632
rect 45836 4072 45888 4078
rect 45836 4014 45888 4020
rect 45560 3664 45612 3670
rect 45560 3606 45612 3612
rect 45652 3664 45704 3670
rect 45652 3606 45704 3612
rect 45192 3460 45244 3466
rect 45192 3402 45244 3408
rect 44916 3120 44968 3126
rect 44916 3062 44968 3068
rect 44548 2576 44600 2582
rect 44548 2518 44600 2524
rect 44456 2372 44508 2378
rect 44456 2314 44508 2320
rect 44560 800 44588 2518
rect 45204 800 45232 3402
rect 45664 2530 45692 3606
rect 45572 2514 45692 2530
rect 45560 2508 45692 2514
rect 45612 2502 45692 2508
rect 45560 2450 45612 2456
rect 45848 800 45876 4014
rect 46492 800 46520 4626
rect 47136 800 47164 5714
rect 47596 5234 47624 7346
rect 47688 6730 47716 7686
rect 47676 6724 47728 6730
rect 47676 6666 47728 6672
rect 49056 6724 49108 6730
rect 49056 6666 49108 6672
rect 48412 6248 48464 6254
rect 48412 6190 48464 6196
rect 47584 5228 47636 5234
rect 47584 5170 47636 5176
rect 47676 5160 47728 5166
rect 47676 5102 47728 5108
rect 47688 2530 47716 5102
rect 47768 3392 47820 3398
rect 47768 3334 47820 3340
rect 47780 2650 47808 3334
rect 47768 2644 47820 2650
rect 47768 2586 47820 2592
rect 47688 2502 47808 2530
rect 47780 800 47808 2502
rect 48424 800 48452 6190
rect 49068 800 49096 6666
rect 726 0 838 800
rect 1370 0 1482 800
rect 2014 0 2126 800
rect 2658 0 2770 800
rect 3302 0 3414 800
rect 3946 0 4058 800
rect 4590 0 4702 800
rect 5234 0 5346 800
rect 5878 0 5990 800
rect 6522 0 6634 800
rect 7166 0 7278 800
rect 7810 0 7922 800
rect 8454 0 8566 800
rect 9098 0 9210 800
rect 9742 0 9854 800
rect 10386 0 10498 800
rect 11030 0 11142 800
rect 11674 0 11786 800
rect 12318 0 12430 800
rect 12962 0 13074 800
rect 13606 0 13718 800
rect 14250 0 14362 800
rect 14894 0 15006 800
rect 15538 0 15650 800
rect 16182 0 16294 800
rect 16826 0 16938 800
rect 17470 0 17582 800
rect 18114 0 18226 800
rect 18758 0 18870 800
rect 19402 0 19514 800
rect 20046 0 20158 800
rect 20690 0 20802 800
rect 21334 0 21446 800
rect 21978 0 22090 800
rect 22622 0 22734 800
rect 23266 0 23378 800
rect 23910 0 24022 800
rect 24554 0 24666 800
rect 25198 0 25310 800
rect 25842 0 25954 800
rect 26486 0 26598 800
rect 27130 0 27242 800
rect 27774 0 27886 800
rect 28418 0 28530 800
rect 29062 0 29174 800
rect 29706 0 29818 800
rect 30350 0 30462 800
rect 30994 0 31106 800
rect 31638 0 31750 800
rect 32282 0 32394 800
rect 32926 0 33038 800
rect 33570 0 33682 800
rect 34214 0 34326 800
rect 34858 0 34970 800
rect 35502 0 35614 800
rect 36146 0 36258 800
rect 36790 0 36902 800
rect 37434 0 37546 800
rect 38078 0 38190 800
rect 38722 0 38834 800
rect 39366 0 39478 800
rect 40010 0 40122 800
rect 40654 0 40766 800
rect 41298 0 41410 800
rect 41942 0 42054 800
rect 42586 0 42698 800
rect 43230 0 43342 800
rect 43874 0 43986 800
rect 44518 0 44630 800
rect 45162 0 45274 800
rect 45806 0 45918 800
rect 46450 0 46562 800
rect 47094 0 47206 800
rect 47738 0 47850 800
rect 48382 0 48494 800
rect 49026 0 49138 800
<< via2 >>
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3054 4120 3110 4176
rect 3698 6296 3754 6352
rect 3974 5616 4030 5672
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4618 5636 4674 5672
rect 4618 5616 4620 5636
rect 4620 5616 4672 5636
rect 4672 5616 4674 5636
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 8114 6296 8170 6352
rect 7010 4120 7066 4176
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
<< metal3 >>
rect 0 47276 800 47516
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 0 45916 800 46156
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 0 44556 800 44796
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 0 43196 800 43436
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 0 41836 800 42076
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 0 40476 800 40716
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 0 39116 800 39356
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 0 37756 800 37996
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 0 36396 800 36636
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 0 35036 800 35276
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 0 33676 800 33916
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 0 32316 800 32556
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 0 30956 800 31196
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 0 29596 800 29836
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 0 28236 800 28476
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 0 26876 800 27116
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 0 25516 800 25756
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 0 24156 800 24396
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 22796 800 23036
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 0 21436 800 21676
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 0 20076 800 20316
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 0 18716 800 18956
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 0 17356 800 17596
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 0 15996 800 16236
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 0 14636 800 14876
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 0 13276 800 13516
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 0 11916 800 12156
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 0 10556 800 10796
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 0 9196 800 9436
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 0 7836 800 8076
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6476 800 6716
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 3693 6354 3759 6357
rect 8109 6354 8175 6357
rect 3693 6352 8175 6354
rect 3693 6296 3698 6352
rect 3754 6296 8114 6352
rect 8170 6296 8175 6352
rect 3693 6294 8175 6296
rect 3693 6291 3759 6294
rect 8109 6291 8175 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 3969 5674 4035 5677
rect 4613 5674 4679 5677
rect 3969 5672 4679 5674
rect 3969 5616 3974 5672
rect 4030 5616 4618 5672
rect 4674 5616 4679 5672
rect 3969 5614 4679 5616
rect 3969 5611 4035 5614
rect 4613 5611 4679 5614
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 0 5116 800 5356
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 3049 4178 3115 4181
rect 7005 4178 7071 4181
rect 3049 4176 7071 4178
rect 3049 4120 3054 4176
rect 3110 4120 7010 4176
rect 7066 4120 7071 4176
rect 3049 4118 7071 4120
rect 3049 4115 3115 4118
rect 7005 4115 7071 4118
rect 0 3756 800 3996
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 0 2396 800 2636
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13248 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1649977179
transform 1 0 9936 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_106 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp 1649977179
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1649977179
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1649977179
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1649977179
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_302
timestamp 1649977179
transform 1 0 28888 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1649977179
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_358
timestamp 1649977179
transform 1 0 34040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_386
timestamp 1649977179
transform 1 0 36616 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_414
timestamp 1649977179
transform 1 0 39192 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_442
timestamp 1649977179
transform 1 0 41768 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_470
timestamp 1649977179
transform 1 0 44344 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_498
timestamp 1649977179
transform 1 0 46920 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_508 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 47840 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_61
timestamp 1649977179
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_83
timestamp 1649977179
transform 1 0 8740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1649977179
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1649977179
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_173
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1649977179
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_229
timestamp 1649977179
transform 1 0 22172 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_251
timestamp 1649977179
transform 1 0 24196 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_302
timestamp 1649977179
transform 1 0 28888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_327
timestamp 1649977179
transform 1 0 31188 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1649977179
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_358
timestamp 1649977179
transform 1 0 34040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_383
timestamp 1649977179
transform 1 0 36340 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1649977179
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_414
timestamp 1649977179
transform 1 0 39192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_439
timestamp 1649977179
transform 1 0 41492 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1649977179
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_470
timestamp 1649977179
transform 1 0 44344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_495
timestamp 1649977179
transform 1 0 46644 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1649977179
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_508
timestamp 1649977179
transform 1 0 47840 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp 1649977179
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1649977179
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_106
timestamp 1649977179
transform 1 0 10856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_131
timestamp 1649977179
transform 1 0 13156 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_163
timestamp 1649977179
transform 1 0 16100 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_218
timestamp 1649977179
transform 1 0 21160 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_222
timestamp 1649977179
transform 1 0 21528 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_244
timestamp 1649977179
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_262
timestamp 1649977179
transform 1 0 25208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_266
timestamp 1649977179
transform 1 0 25576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_288
timestamp 1649977179
transform 1 0 27600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_295
timestamp 1649977179
transform 1 0 28244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_302
timestamp 1649977179
transform 1 0 28888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_330
timestamp 1649977179
transform 1 0 31464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_355
timestamp 1649977179
transform 1 0 33764 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1649977179
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_386
timestamp 1649977179
transform 1 0 36616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_411
timestamp 1649977179
transform 1 0 38916 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_442
timestamp 1649977179
transform 1 0 41768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_467
timestamp 1649977179
transform 1 0 44068 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1649977179
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_498
timestamp 1649977179
transform 1 0 46920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_505
timestamp 1649977179
transform 1 0 47564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1649977179
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_26
timestamp 1649977179
transform 1 0 3496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_30
timestamp 1649977179
transform 1 0 3864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_61
timestamp 1649977179
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_83
timestamp 1649977179
transform 1 0 8740 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_117
timestamp 1649977179
transform 1 0 11868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_128
timestamp 1649977179
transform 1 0 12880 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_153
timestamp 1649977179
transform 1 0 15180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_178
timestamp 1649977179
transform 1 0 17480 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_185
timestamp 1649977179
transform 1 0 18124 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_210
timestamp 1649977179
transform 1 0 20424 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1649977179
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_228
timestamp 1649977179
transform 1 0 22080 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_235
timestamp 1649977179
transform 1 0 22724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1649977179
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_268
timestamp 1649977179
transform 1 0 25760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_275
timestamp 1649977179
transform 1 0 26404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_284
timestamp 1649977179
transform 1 0 27232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_291
timestamp 1649977179
transform 1 0 27876 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_316
timestamp 1649977179
transform 1 0 30176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_323
timestamp 1649977179
transform 1 0 30820 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1649977179
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_358
timestamp 1649977179
transform 1 0 34040 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_364
timestamp 1649977179
transform 1 0 34592 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_386
timestamp 1649977179
transform 1 0 36616 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_415
timestamp 1649977179
transform 1 0 39284 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_444
timestamp 1649977179
transform 1 0 41952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_472
timestamp 1649977179
transform 1 0 44528 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_476
timestamp 1649977179
transform 1 0 44896 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_498
timestamp 1649977179
transform 1 0 46920 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_508
timestamp 1649977179
transform 1 0 47840 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_8
timestamp 1649977179
transform 1 0 1840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_50
timestamp 1649977179
transform 1 0 5704 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_106
timestamp 1649977179
transform 1 0 10856 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1649977179
transform 1 0 14812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_157
timestamp 1649977179
transform 1 0 15548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_164
timestamp 1649977179
transform 1 0 16192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_171
timestamp 1649977179
transform 1 0 16836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_178
timestamp 1649977179
transform 1 0 17480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_185
timestamp 1649977179
transform 1 0 18124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1649977179
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_204
timestamp 1649977179
transform 1 0 19872 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_218
timestamp 1649977179
transform 1 0 21160 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_227
timestamp 1649977179
transform 1 0 21988 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_234
timestamp 1649977179
transform 1 0 22632 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_241
timestamp 1649977179
transform 1 0 23276 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1649977179
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_258
timestamp 1649977179
transform 1 0 24840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_272
timestamp 1649977179
transform 1 0 26128 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_280
timestamp 1649977179
transform 1 0 26864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_286
timestamp 1649977179
transform 1 0 27416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_294
timestamp 1649977179
transform 1 0 28152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_312
timestamp 1649977179
transform 1 0 29808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_319
timestamp 1649977179
transform 1 0 30452 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_326
timestamp 1649977179
transform 1 0 31096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_334
timestamp 1649977179
transform 1 0 31832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_339
timestamp 1649977179
transform 1 0 32292 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_351
timestamp 1649977179
transform 1 0 33396 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_358
timestamp 1649977179
transform 1 0 34040 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_368
timestamp 1649977179
transform 1 0 34960 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_375
timestamp 1649977179
transform 1 0 35604 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_382
timestamp 1649977179
transform 1 0 36248 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_399
timestamp 1649977179
transform 1 0 37812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_406
timestamp 1649977179
transform 1 0 38456 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_424
timestamp 1649977179
transform 1 0 40112 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_434
timestamp 1649977179
transform 1 0 41032 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_441
timestamp 1649977179
transform 1 0 41676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_448
timestamp 1649977179
transform 1 0 42320 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_455
timestamp 1649977179
transform 1 0 42964 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_462
timestamp 1649977179
transform 1 0 43608 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_472
timestamp 1649977179
transform 1 0 44528 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_482
timestamp 1649977179
transform 1 0 45448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_507
timestamp 1649977179
transform 1 0 47748 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_515
timestamp 1649977179
transform 1 0 48484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_19
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1649977179
transform 1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp 1649977179
transform 1 0 3864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_41
timestamp 1649977179
transform 1 0 4876 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_61
timestamp 1649977179
transform 1 0 6716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_97
timestamp 1649977179
transform 1 0 10028 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_133
timestamp 1649977179
transform 1 0 13340 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_141
timestamp 1649977179
transform 1 0 14076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 1649977179
transform 1 0 14444 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_153
timestamp 1649977179
transform 1 0 15180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_160
timestamp 1649977179
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_172
timestamp 1649977179
transform 1 0 16928 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_179
timestamp 1649977179
transform 1 0 17572 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_190
timestamp 1649977179
transform 1 0 18584 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1649977179
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_204
timestamp 1649977179
transform 1 0 19872 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_211
timestamp 1649977179
transform 1 0 20516 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1649977179
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_228
timestamp 1649977179
transform 1 0 22080 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1649977179
transform 1 0 22816 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_241
timestamp 1649977179
transform 1 0 23276 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1649977179
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_251
timestamp 1649977179
transform 1 0 24196 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_258 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24840 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_270
timestamp 1649977179
transform 1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1649977179
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_299
timestamp 1649977179
transform 1 0 28612 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_306
timestamp 1649977179
transform 1 0 29256 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_318
timestamp 1649977179
transform 1 0 30360 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_322
timestamp 1649977179
transform 1 0 30728 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_340
timestamp 1649977179
transform 1 0 32384 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_347
timestamp 1649977179
transform 1 0 33028 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_354
timestamp 1649977179
transform 1 0 33672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_368
timestamp 1649977179
transform 1 0 34960 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_375
timestamp 1649977179
transform 1 0 35604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_382
timestamp 1649977179
transform 1 0 36248 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp 1649977179
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_396
timestamp 1649977179
transform 1 0 37536 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1649977179
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_410
timestamp 1649977179
transform 1 0 38824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_424
timestamp 1649977179
transform 1 0 40112 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_431
timestamp 1649977179
transform 1 0 40756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_438
timestamp 1649977179
transform 1 0 41400 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_446
timestamp 1649977179
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_452
timestamp 1649977179
transform 1 0 42688 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_459
timestamp 1649977179
transform 1 0 43332 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_466
timestamp 1649977179
transform 1 0 43976 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1649977179
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_508
timestamp 1649977179
transform 1 0 47840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_10
timestamp 1649977179
transform 1 0 2024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_17
timestamp 1649977179
transform 1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1649977179
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1649977179
transform 1 0 4048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_56
timestamp 1649977179
transform 1 0 6256 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_92
timestamp 1649977179
transform 1 0 9568 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_100
timestamp 1649977179
transform 1 0 10304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_108
timestamp 1649977179
transform 1 0 11040 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_117
timestamp 1649977179
transform 1 0 11868 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_125
timestamp 1649977179
transform 1 0 12604 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_146
timestamp 1649977179
transform 1 0 14536 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_326
timestamp 1649977179
transform 1 0 31096 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_340
timestamp 1649977179
transform 1 0 32384 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_352
timestamp 1649977179
transform 1 0 33488 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_384
timestamp 1649977179
transform 1 0 36432 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_391
timestamp 1649977179
transform 1 0 37076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_406
timestamp 1649977179
transform 1 0 38456 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_418
timestamp 1649977179
transform 1 0 39560 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_426
timestamp 1649977179
transform 1 0 40296 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_441
timestamp 1649977179
transform 1 0 41676 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_453
timestamp 1649977179
transform 1 0 42780 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_462
timestamp 1649977179
transform 1 0 43608 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_468
timestamp 1649977179
transform 1 0 44160 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_472
timestamp 1649977179
transform 1 0 44528 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_480
timestamp 1649977179
transform 1 0 45264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_487
timestamp 1649977179
transform 1 0 45908 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_512
timestamp 1649977179
transform 1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_12
timestamp 1649977179
transform 1 0 2208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_19
timestamp 1649977179
transform 1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_26
timestamp 1649977179
transform 1 0 3496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_33
timestamp 1649977179
transform 1 0 4140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_40
timestamp 1649977179
transform 1 0 4784 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_49
timestamp 1649977179
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_77
timestamp 1649977179
transform 1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_84
timestamp 1649977179
transform 1 0 8832 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_94
timestamp 1649977179
transform 1 0 9752 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_140
timestamp 1649977179
transform 1 0 13984 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_147
timestamp 1649977179
transform 1 0 14628 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_159
timestamp 1649977179
transform 1 0 15732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1649977179
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1649977179
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1649977179
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_500
timestamp 1649977179
transform 1 0 47104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_508
timestamp 1649977179
transform 1 0 47840 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_12
timestamp 1649977179
transform 1 0 2208 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_20
timestamp 1649977179
transform 1 0 2944 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1649977179
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_33
timestamp 1649977179
transform 1 0 4140 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_40
timestamp 1649977179
transform 1 0 4784 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_64
timestamp 1649977179
transform 1 0 6992 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 1649977179
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1649977179
transform 1 0 9200 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_95
timestamp 1649977179
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_99
timestamp 1649977179
transform 1 0 10212 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_120
timestamp 1649977179
transform 1 0 12144 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_128
timestamp 1649977179
transform 1 0 12880 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1649977179
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1649977179
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1649977179
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1649977179
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1649977179
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_12
timestamp 1649977179
transform 1 0 2208 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_20
timestamp 1649977179
transform 1 0 2944 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_25
timestamp 1649977179
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_37
timestamp 1649977179
transform 1 0 4508 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_41
timestamp 1649977179
transform 1 0 4876 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 1649977179
transform 1 0 5244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1649977179
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_73
timestamp 1649977179
transform 1 0 7820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_94
timestamp 1649977179
transform 1 0 9752 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_102
timestamp 1649977179
transform 1 0 10488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp 1649977179
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_116
timestamp 1649977179
transform 1 0 11776 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_128
timestamp 1649977179
transform 1 0 12880 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_140
timestamp 1649977179
transform 1 0 13984 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_152
timestamp 1649977179
transform 1 0 15088 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1649977179
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1649977179
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1649977179
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1649977179
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_489
timestamp 1649977179
transform 1 0 46092 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_493
timestamp 1649977179
transform 1 0 46460 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_500
timestamp 1649977179
transform 1 0 47104 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_508
timestamp 1649977179
transform 1 0 47840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_9
timestamp 1649977179
transform 1 0 1932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_13
timestamp 1649977179
transform 1 0 2300 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_17
timestamp 1649977179
transform 1 0 2668 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1649977179
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_57
timestamp 1649977179
transform 1 0 6348 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_63
timestamp 1649977179
transform 1 0 6900 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_67
timestamp 1649977179
transform 1 0 7268 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_75
timestamp 1649977179
transform 1 0 8004 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp 1649977179
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_93
timestamp 1649977179
transform 1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_98
timestamp 1649977179
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_103
timestamp 1649977179
transform 1 0 10580 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_110
timestamp 1649977179
transform 1 0 11224 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_122
timestamp 1649977179
transform 1 0 12328 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1649977179
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1649977179
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1649977179
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_497
timestamp 1649977179
transform 1 0 46828 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_508
timestamp 1649977179
transform 1 0 47840 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_9
timestamp 1649977179
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_21
timestamp 1649977179
transform 1 0 3036 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_33
timestamp 1649977179
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_45
timestamp 1649977179
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1649977179
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_74
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_78
timestamp 1649977179
transform 1 0 8280 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_82
timestamp 1649977179
transform 1 0 8648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_89
timestamp 1649977179
transform 1 0 9292 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_96
timestamp 1649977179
transform 1 0 9936 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1649977179
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1649977179
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1649977179
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1649977179
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_511
timestamp 1649977179
transform 1 0 48116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_515
timestamp 1649977179
transform 1 0 48484 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_103
timestamp 1649977179
transform 1 0 10580 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_115
timestamp 1649977179
transform 1 0 11684 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_123
timestamp 1649977179
transform 1 0 12420 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_127
timestamp 1649977179
transform 1 0 12788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1649977179
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1649977179
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1649977179
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1649977179
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1649977179
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1649977179
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1649977179
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1649977179
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1649977179
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1649977179
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1649977179
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1649977179
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1649977179
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1649977179
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1649977179
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_513
timestamp 1649977179
transform 1 0 48300 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1649977179
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1649977179
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1649977179
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1649977179
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1649977179
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1649977179
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1649977179
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1649977179
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1649977179
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_513
timestamp 1649977179
transform 1 0 48300 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1649977179
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1649977179
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1649977179
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1649977179
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1649977179
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1649977179
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1649977179
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1649977179
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1649977179
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1649977179
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1649977179
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1649977179
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1649977179
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1649977179
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1649977179
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1649977179
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1649977179
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1649977179
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1649977179
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_513
timestamp 1649977179
transform 1 0 48300 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1649977179
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1649977179
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1649977179
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1649977179
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1649977179
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1649977179
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1649977179
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1649977179
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1649977179
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1649977179
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1649977179
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_513
timestamp 1649977179
transform 1 0 48300 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1649977179
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1649977179
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1649977179
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1649977179
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1649977179
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1649977179
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1649977179
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1649977179
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1649977179
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_513
timestamp 1649977179
transform 1 0 48300 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1649977179
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1649977179
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1649977179
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1649977179
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1649977179
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1649977179
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1649977179
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1649977179
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1649977179
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1649977179
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1649977179
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_513
timestamp 1649977179
transform 1 0 48300 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1649977179
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1649977179
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1649977179
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1649977179
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1649977179
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1649977179
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1649977179
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1649977179
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1649977179
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1649977179
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1649977179
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1649977179
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1649977179
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_513
timestamp 1649977179
transform 1 0 48300 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1649977179
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1649977179
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1649977179
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1649977179
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1649977179
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1649977179
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1649977179
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1649977179
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1649977179
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1649977179
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1649977179
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1649977179
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1649977179
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1649977179
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1649977179
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1649977179
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_513
timestamp 1649977179
transform 1 0 48300 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1649977179
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1649977179
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1649977179
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1649977179
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1649977179
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1649977179
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1649977179
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1649977179
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1649977179
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1649977179
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1649977179
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1649977179
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1649977179
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1649977179
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1649977179
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1649977179
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_513
timestamp 1649977179
transform 1 0 48300 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1649977179
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1649977179
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1649977179
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1649977179
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1649977179
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1649977179
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1649977179
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1649977179
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1649977179
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1649977179
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1649977179
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1649977179
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1649977179
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_513
timestamp 1649977179
transform 1 0 48300 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1649977179
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1649977179
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1649977179
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1649977179
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1649977179
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1649977179
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1649977179
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1649977179
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1649977179
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1649977179
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1649977179
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1649977179
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1649977179
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_513
timestamp 1649977179
transform 1 0 48300 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1649977179
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1649977179
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1649977179
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1649977179
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1649977179
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1649977179
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1649977179
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1649977179
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1649977179
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1649977179
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1649977179
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1649977179
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1649977179
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1649977179
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1649977179
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1649977179
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1649977179
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1649977179
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1649977179
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_513
timestamp 1649977179
transform 1 0 48300 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1649977179
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1649977179
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1649977179
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1649977179
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1649977179
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1649977179
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1649977179
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1649977179
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1649977179
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1649977179
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1649977179
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1649977179
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1649977179
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1649977179
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1649977179
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1649977179
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1649977179
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1649977179
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1649977179
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1649977179
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1649977179
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1649977179
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1649977179
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1649977179
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1649977179
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1649977179
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1649977179
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1649977179
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1649977179
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_513
timestamp 1649977179
transform 1 0 48300 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1649977179
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1649977179
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1649977179
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1649977179
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1649977179
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1649977179
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1649977179
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1649977179
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1649977179
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1649977179
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1649977179
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1649977179
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1649977179
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1649977179
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1649977179
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1649977179
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1649977179
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_513
timestamp 1649977179
transform 1 0 48300 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1649977179
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1649977179
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1649977179
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1649977179
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1649977179
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1649977179
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1649977179
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1649977179
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1649977179
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1649977179
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1649977179
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1649977179
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1649977179
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1649977179
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1649977179
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1649977179
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1649977179
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1649977179
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1649977179
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1649977179
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1649977179
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1649977179
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1649977179
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1649977179
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1649977179
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1649977179
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1649977179
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1649977179
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1649977179
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1649977179
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1649977179
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1649977179
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1649977179
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1649977179
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1649977179
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1649977179
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1649977179
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1649977179
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1649977179
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1649977179
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1649977179
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1649977179
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1649977179
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1649977179
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1649977179
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1649977179
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1649977179
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1649977179
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1649977179
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1649977179
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1649977179
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1649977179
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1649977179
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1649977179
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1649977179
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1649977179
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1649977179
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1649977179
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1649977179
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1649977179
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1649977179
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1649977179
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1649977179
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1649977179
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1649977179
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_513
timestamp 1649977179
transform 1 0 48300 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1649977179
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1649977179
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1649977179
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1649977179
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1649977179
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1649977179
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1649977179
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1649977179
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1649977179
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1649977179
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1649977179
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1649977179
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1649977179
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1649977179
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1649977179
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1649977179
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1649977179
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1649977179
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1649977179
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1649977179
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1649977179
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1649977179
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1649977179
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1649977179
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1649977179
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1649977179
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1649977179
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1649977179
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1649977179
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1649977179
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1649977179
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1649977179
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1649977179
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1649977179
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1649977179
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1649977179
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1649977179
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1649977179
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1649977179
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1649977179
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1649977179
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1649977179
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1649977179
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1649977179
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1649977179
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1649977179
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_513
timestamp 1649977179
transform 1 0 48300 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1649977179
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1649977179
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1649977179
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1649977179
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1649977179
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1649977179
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1649977179
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1649977179
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1649977179
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1649977179
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1649977179
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1649977179
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1649977179
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1649977179
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1649977179
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1649977179
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1649977179
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1649977179
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1649977179
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1649977179
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1649977179
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1649977179
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1649977179
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1649977179
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1649977179
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1649977179
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1649977179
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1649977179
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1649977179
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1649977179
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1649977179
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1649977179
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1649977179
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1649977179
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1649977179
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1649977179
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1649977179
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1649977179
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1649977179
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1649977179
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1649977179
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1649977179
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1649977179
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1649977179
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1649977179
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1649977179
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1649977179
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1649977179
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1649977179
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1649977179
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1649977179
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1649977179
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1649977179
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1649977179
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1649977179
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1649977179
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1649977179
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1649977179
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1649977179
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1649977179
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1649977179
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1649977179
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1649977179
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1649977179
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1649977179
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1649977179
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1649977179
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1649977179
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1649977179
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1649977179
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1649977179
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1649977179
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1649977179
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1649977179
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1649977179
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1649977179
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1649977179
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1649977179
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1649977179
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_513
timestamp 1649977179
transform 1 0 48300 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1649977179
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1649977179
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1649977179
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1649977179
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1649977179
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1649977179
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1649977179
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1649977179
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1649977179
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1649977179
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1649977179
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1649977179
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1649977179
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1649977179
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1649977179
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1649977179
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1649977179
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1649977179
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1649977179
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1649977179
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_513
timestamp 1649977179
transform 1 0 48300 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1649977179
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1649977179
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1649977179
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1649977179
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1649977179
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1649977179
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1649977179
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1649977179
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1649977179
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1649977179
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1649977179
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1649977179
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1649977179
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1649977179
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1649977179
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1649977179
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1649977179
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1649977179
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1649977179
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1649977179
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_513
timestamp 1649977179
transform 1 0 48300 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1649977179
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1649977179
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1649977179
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1649977179
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1649977179
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1649977179
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1649977179
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1649977179
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1649977179
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1649977179
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1649977179
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1649977179
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1649977179
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1649977179
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_513
timestamp 1649977179
transform 1 0 48300 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1649977179
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1649977179
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1649977179
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1649977179
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1649977179
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1649977179
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1649977179
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1649977179
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1649977179
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1649977179
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1649977179
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1649977179
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1649977179
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1649977179
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_513
timestamp 1649977179
transform 1 0 48300 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1649977179
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1649977179
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1649977179
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1649977179
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1649977179
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1649977179
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1649977179
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1649977179
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1649977179
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1649977179
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1649977179
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1649977179
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1649977179
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1649977179
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1649977179
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1649977179
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1649977179
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1649977179
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1649977179
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_513
timestamp 1649977179
transform 1 0 48300 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1649977179
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1649977179
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1649977179
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1649977179
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1649977179
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1649977179
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1649977179
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1649977179
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1649977179
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1649977179
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1649977179
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1649977179
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1649977179
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1649977179
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_513
timestamp 1649977179
transform 1 0 48300 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1649977179
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1649977179
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1649977179
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1649977179
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1649977179
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1649977179
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1649977179
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1649977179
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1649977179
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1649977179
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1649977179
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1649977179
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1649977179
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1649977179
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1649977179
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1649977179
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1649977179
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1649977179
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1649977179
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1649977179
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_513
timestamp 1649977179
transform 1 0 48300 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1649977179
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1649977179
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1649977179
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1649977179
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1649977179
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1649977179
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1649977179
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1649977179
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1649977179
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1649977179
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1649977179
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1649977179
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1649977179
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1649977179
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1649977179
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1649977179
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1649977179
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1649977179
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1649977179
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1649977179
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1649977179
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1649977179
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1649977179
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1649977179
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1649977179
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1649977179
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1649977179
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1649977179
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1649977179
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1649977179
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1649977179
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1649977179
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_513
timestamp 1649977179
transform 1 0 48300 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1649977179
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1649977179
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1649977179
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1649977179
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1649977179
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1649977179
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1649977179
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1649977179
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1649977179
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1649977179
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1649977179
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1649977179
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1649977179
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1649977179
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1649977179
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1649977179
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1649977179
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1649977179
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1649977179
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1649977179
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1649977179
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1649977179
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1649977179
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1649977179
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1649977179
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1649977179
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1649977179
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1649977179
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1649977179
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1649977179
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1649977179
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1649977179
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1649977179
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1649977179
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1649977179
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1649977179
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1649977179
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1649977179
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1649977179
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_513
timestamp 1649977179
transform 1 0 48300 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1649977179
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1649977179
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1649977179
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1649977179
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1649977179
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1649977179
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1649977179
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1649977179
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1649977179
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1649977179
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1649977179
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1649977179
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1649977179
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1649977179
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1649977179
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1649977179
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1649977179
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1649977179
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1649977179
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1649977179
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1649977179
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1649977179
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1649977179
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1649977179
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1649977179
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1649977179
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1649977179
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1649977179
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1649977179
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1649977179
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1649977179
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1649977179
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1649977179
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1649977179
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1649977179
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1649977179
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_513
timestamp 1649977179
transform 1 0 48300 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1649977179
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1649977179
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1649977179
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1649977179
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1649977179
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1649977179
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1649977179
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1649977179
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1649977179
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1649977179
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1649977179
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1649977179
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1649977179
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1649977179
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1649977179
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1649977179
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1649977179
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1649977179
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1649977179
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1649977179
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1649977179
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1649977179
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1649977179
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1649977179
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1649977179
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1649977179
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1649977179
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1649977179
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1649977179
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1649977179
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1649977179
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1649977179
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1649977179
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1649977179
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1649977179
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1649977179
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1649977179
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1649977179
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1649977179
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_513
timestamp 1649977179
transform 1 0 48300 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1649977179
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1649977179
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1649977179
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1649977179
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1649977179
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1649977179
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1649977179
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1649977179
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1649977179
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1649977179
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1649977179
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1649977179
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1649977179
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1649977179
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1649977179
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1649977179
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1649977179
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1649977179
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1649977179
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1649977179
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1649977179
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1649977179
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1649977179
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1649977179
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1649977179
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1649977179
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1649977179
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1649977179
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1649977179
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1649977179
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1649977179
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1649977179
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1649977179
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1649977179
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1649977179
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1649977179
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1649977179
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1649977179
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1649977179
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1649977179
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1649977179
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1649977179
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1649977179
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1649977179
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1649977179
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1649977179
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1649977179
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1649977179
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1649977179
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1649977179
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1649977179
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1649977179
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1649977179
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1649977179
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1649977179
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1649977179
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1649977179
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1649977179
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1649977179
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1649977179
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1649977179
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1649977179
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1649977179
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1649977179
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1649977179
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1649977179
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1649977179
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1649977179
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1649977179
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1649977179
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1649977179
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1649977179
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_513
timestamp 1649977179
transform 1 0 48300 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1649977179
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1649977179
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1649977179
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1649977179
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1649977179
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1649977179
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1649977179
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1649977179
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1649977179
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1649977179
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1649977179
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1649977179
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1649977179
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1649977179
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1649977179
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1649977179
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1649977179
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1649977179
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1649977179
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1649977179
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1649977179
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1649977179
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1649977179
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1649977179
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1649977179
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1649977179
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1649977179
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1649977179
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1649977179
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1649977179
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1649977179
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1649977179
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1649977179
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1649977179
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1649977179
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1649977179
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1649977179
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_513
timestamp 1649977179
transform 1 0 48300 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1649977179
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1649977179
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1649977179
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1649977179
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1649977179
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1649977179
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1649977179
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1649977179
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1649977179
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1649977179
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1649977179
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1649977179
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1649977179
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1649977179
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1649977179
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1649977179
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1649977179
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1649977179
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1649977179
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1649977179
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1649977179
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1649977179
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1649977179
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1649977179
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1649977179
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1649977179
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1649977179
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1649977179
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1649977179
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1649977179
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1649977179
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1649977179
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1649977179
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1649977179
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1649977179
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_513
timestamp 1649977179
transform 1 0 48300 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1649977179
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1649977179
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1649977179
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1649977179
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1649977179
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1649977179
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1649977179
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1649977179
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1649977179
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1649977179
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1649977179
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1649977179
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1649977179
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1649977179
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1649977179
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1649977179
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1649977179
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1649977179
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1649977179
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1649977179
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1649977179
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1649977179
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1649977179
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1649977179
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1649977179
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1649977179
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1649977179
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1649977179
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1649977179
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1649977179
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1649977179
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1649977179
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1649977179
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1649977179
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1649977179
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1649977179
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1649977179
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1649977179
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1649977179
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1649977179
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1649977179
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1649977179
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1649977179
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1649977179
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1649977179
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1649977179
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1649977179
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1649977179
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_513
timestamp 1649977179
transform 1 0 48300 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1649977179
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1649977179
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1649977179
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1649977179
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1649977179
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1649977179
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1649977179
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1649977179
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1649977179
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1649977179
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1649977179
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1649977179
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1649977179
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1649977179
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1649977179
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1649977179
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_513
timestamp 1649977179
transform 1 0 48300 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1649977179
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1649977179
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1649977179
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1649977179
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1649977179
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1649977179
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1649977179
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1649977179
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1649977179
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1649977179
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1649977179
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1649977179
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1649977179
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1649977179
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_513
timestamp 1649977179
transform 1 0 48300 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1649977179
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1649977179
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1649977179
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1649977179
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1649977179
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1649977179
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1649977179
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1649977179
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_513
timestamp 1649977179
transform 1 0 48300 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1649977179
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1649977179
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1649977179
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1649977179
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1649977179
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1649977179
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1649977179
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1649977179
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1649977179
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1649977179
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1649977179
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1649977179
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1649977179
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1649977179
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1649977179
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1649977179
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_513
timestamp 1649977179
transform 1 0 48300 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1649977179
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1649977179
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1649977179
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1649977179
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1649977179
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1649977179
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1649977179
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1649977179
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1649977179
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1649977179
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1649977179
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1649977179
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1649977179
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1649977179
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1649977179
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1649977179
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1649977179
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1649977179
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1649977179
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_513
timestamp 1649977179
transform 1 0 48300 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1649977179
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1649977179
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1649977179
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1649977179
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1649977179
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1649977179
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1649977179
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1649977179
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1649977179
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1649977179
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1649977179
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1649977179
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1649977179
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1649977179
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1649977179
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1649977179
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1649977179
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1649977179
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1649977179
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1649977179
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1649977179
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1649977179
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1649977179
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1649977179
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1649977179
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1649977179
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1649977179
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_505
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_513
timestamp 1649977179
transform 1 0 48300 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1649977179
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1649977179
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1649977179
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1649977179
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1649977179
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1649977179
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1649977179
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1649977179
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1649977179
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1649977179
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1649977179
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1649977179
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1649977179
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1649977179
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1649977179
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1649977179
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1649977179
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1649977179
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1649977179
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1649977179
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1649977179
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1649977179
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1649977179
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1649977179
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1649977179
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1649977179
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1649977179
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1649977179
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1649977179
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_513
timestamp 1649977179
transform 1 0 48300 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1649977179
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1649977179
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1649977179
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1649977179
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1649977179
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1649977179
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1649977179
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1649977179
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1649977179
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1649977179
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1649977179
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1649977179
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1649977179
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1649977179
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1649977179
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1649977179
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1649977179
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1649977179
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1649977179
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1649977179
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1649977179
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1649977179
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1649977179
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1649977179
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1649977179
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1649977179
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1649977179
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1649977179
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1649977179
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1649977179
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1649977179
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1649977179
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_505
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_513
timestamp 1649977179
transform 1 0 48300 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_3
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_7
timestamp 1649977179
transform 1 0 1748 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_12
timestamp 1649977179
transform 1 0 2208 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_24
timestamp 1649977179
transform 1 0 3312 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_82_50
timestamp 1649977179
transform 1 0 5704 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_82_57
timestamp 1649977179
transform 1 0 6348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_69
timestamp 1649977179
transform 1 0 7452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_81
timestamp 1649977179
transform 1 0 8556 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1649977179
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_109
timestamp 1649977179
transform 1 0 11132 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_113
timestamp 1649977179
transform 1 0 11500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_125
timestamp 1649977179
transform 1 0 12604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1649977179
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_165
timestamp 1649977179
transform 1 0 16284 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_169
timestamp 1649977179
transform 1 0 16652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_181
timestamp 1649977179
transform 1 0 17756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_193
timestamp 1649977179
transform 1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_229
timestamp 1649977179
transform 1 0 22172 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_241
timestamp 1649977179
transform 1 0 23276 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_249
timestamp 1649977179
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_82_253
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_259
timestamp 1649977179
transform 1 0 24932 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_264
timestamp 1649977179
transform 1 0 25392 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_276
timestamp 1649977179
transform 1 0 26496 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_281
timestamp 1649977179
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_293
timestamp 1649977179
transform 1 0 28060 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_300
timestamp 1649977179
transform 1 0 28704 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1649977179
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_333
timestamp 1649977179
transform 1 0 31740 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_341
timestamp 1649977179
transform 1 0 32476 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_353
timestamp 1649977179
transform 1 0 33580 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1649977179
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_372
timestamp 1649977179
transform 1 0 35328 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_384
timestamp 1649977179
transform 1 0 36432 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_82_393
timestamp 1649977179
transform 1 0 37260 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_401
timestamp 1649977179
transform 1 0 37996 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_408
timestamp 1649977179
transform 1 0 38640 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_449
timestamp 1649977179
transform 1 0 42412 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_459
timestamp 1649977179
transform 1 0 43332 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_471
timestamp 1649977179
transform 1 0 44436 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1649977179
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_487
timestamp 1649977179
transform 1 0 45908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_499
timestamp 1649977179
transform 1 0 47012 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_503
timestamp 1649977179
transform 1 0 47380 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_505
timestamp 1649977179
transform 1 0 47564 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_512
timestamp 1649977179
transform 1 0 48208 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 42320 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 47472 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _180_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19504 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1649977179
transform 1 0 44160 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 47564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1649977179
transform 1 0 47840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1649977179
transform 1 0 45632 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _187_
timestamp 1649977179
transform 1 0 45080 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1649977179
transform 1 0 47932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1649977179
transform 1 0 44344 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1649977179
transform 1 0 43332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1649977179
transform 1 0 43700 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _193_
timestamp 1649977179
transform 1 0 40664 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _194_
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _195_
timestamp 1649977179
transform 1 0 42688 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1649977179
transform 1 0 41124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _197_
timestamp 1649977179
transform 1 0 41400 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _198_
timestamp 1649977179
transform 1 0 40480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _199_
timestamp 1649977179
transform 1 0 37444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1649977179
transform 1 0 38548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 1649977179
transform 1 0 37904 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1649977179
transform 1 0 38180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20240 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _206_
timestamp 1649977179
transform 1 0 33028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _207_
timestamp 1649977179
transform 1 0 36616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _208_
timestamp 1649977179
transform 1 0 35328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _209_
timestamp 1649977179
transform 1 0 35328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _210_
timestamp 1649977179
transform 1 0 34040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1649977179
transform 1 0 33396 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _212_
timestamp 1649977179
transform 1 0 31924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _213_
timestamp 1649977179
transform 1 0 32752 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1649977179
transform 1 0 31096 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1649977179
transform 1 0 30452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1649977179
transform 1 0 31188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _218_
timestamp 1649977179
transform 1 0 27784 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1649977179
transform 1 0 28980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1649977179
transform 1 0 28336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1649977179
transform 1 0 28520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1649977179
transform 1 0 27600 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1649977179
transform 1 0 27968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _224_
timestamp 1649977179
transform 1 0 23092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1649977179
transform 1 0 25208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1649977179
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1649977179
transform 1 0 22448 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1649977179
transform 1 0 23000 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _230_
timestamp 1649977179
transform 1 0 20792 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1649977179
transform 1 0 22356 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1649977179
transform 1 0 20240 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1649977179
transform 1 0 17848 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _236_
timestamp 1649977179
transform -1 0 12880 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _237_
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1649977179
transform 1 0 17204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1649977179
transform 1 0 17296 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1649977179
transform 1 0 15272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _243_
timestamp 1649977179
transform 1 0 14444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1649977179
transform 1 0 14260 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1649977179
transform 1 0 14352 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1649977179
transform 1 0 14904 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _249_
timestamp 1649977179
transform 1 0 12236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1649977179
transform 1 0 10672 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1649977179
transform 1 0 10948 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _255_
timestamp 1649977179
transform 1 0 12972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1649977179
transform 1 0 9384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1649977179
transform 1 0 8372 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1649977179
transform 1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1649977179
transform 1 0 2944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1649977179
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1649977179
transform 1 0 6072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1649977179
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1649977179
transform 1 0 3864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1649977179
transform 1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _267_
timestamp 1649977179
transform 1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1649977179
transform 1 0 2576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1649977179
transform 1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1649977179
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1649977179
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1649977179
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1649977179
transform 1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1649977179
transform 1 0 4968 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5152 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4232 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6808 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5244 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7544 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _283_
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11408 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9384 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _288_
timestamp 1649977179
transform 1 0 10120 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _289_
timestamp 1649977179
transform 1 0 10120 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _290_
timestamp 1649977179
transform 1 0 10396 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _291_
timestamp 1649977179
transform 1 0 8096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1649977179
transform 1 0 6992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1649977179
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1649977179
transform 1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1649977179
transform 1 0 10304 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1649977179
transform 1 0 12512 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1649977179
transform 1 0 13064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _300_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5152 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _301_
timestamp 1649977179
transform 1 0 4416 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _302_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _303_
timestamp 1649977179
transform 1 0 6624 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _304_
timestamp 1649977179
transform 1 0 7820 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _305_
timestamp 1649977179
transform 1 0 7912 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _306_
timestamp 1649977179
transform 1 0 10304 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _307_
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  _368_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9108 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _369_
timestamp 1649977179
transform 1 0 9108 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _370_
timestamp 1649977179
transform 1 0 11224 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _371_
timestamp 1649977179
transform 1 0 11408 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _372_
timestamp 1649977179
transform 1 0 11592 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _373_
timestamp 1649977179
transform 1 0 11960 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _374_
timestamp 1649977179
transform 1 0 13248 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _375__15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14168 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _375_
timestamp 1649977179
transform 1 0 14168 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _376__16
timestamp 1649977179
transform 1 0 14904 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _376_
timestamp 1649977179
transform 1 0 14260 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _377__17
timestamp 1649977179
transform 1 0 15548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _377_
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _378__18
timestamp 1649977179
transform 1 0 15916 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _378_
timestamp 1649977179
transform 1 0 16468 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _379__19
timestamp 1649977179
transform 1 0 16560 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _379_
timestamp 1649977179
transform 1 0 16836 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _380__20
timestamp 1649977179
transform 1 0 17204 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _380_
timestamp 1649977179
transform 1 0 17112 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _381__21
timestamp 1649977179
transform 1 0 17848 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _381_
timestamp 1649977179
transform 1 0 18492 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _382__22
timestamp 1649977179
transform 1 0 18952 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _382_
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _383__23
timestamp 1649977179
transform 1 0 19596 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _383_
timestamp 1649977179
transform 1 0 19412 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _384__24
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _384_
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _385__25
timestamp 1649977179
transform 1 0 21712 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _385_
timestamp 1649977179
transform 1 0 21620 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _386__26
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _386_
timestamp 1649977179
transform 1 0 21988 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _387__27
timestamp 1649977179
transform 1 0 23000 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _387_
timestamp 1649977179
transform 1 0 22264 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _388__28
timestamp 1649977179
transform 1 0 23920 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _388_
timestamp 1649977179
transform 1 0 23828 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _389__29
timestamp 1649977179
transform 1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _389_
timestamp 1649977179
transform 1 0 24564 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _390__30
timestamp 1649977179
transform 1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _390_
timestamp 1649977179
transform 1 0 24564 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _391__31
timestamp 1649977179
transform 1 0 26128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _391_
timestamp 1649977179
transform 1 0 25668 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _392__32
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _392_
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _393__33
timestamp 1649977179
transform 1 0 28612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _393_
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _394__34
timestamp 1649977179
transform 1 0 27140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _394_
timestamp 1649977179
transform 1 0 29256 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _395__35
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _395_
timestamp 1649977179
transform 1 0 28244 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _396__36
timestamp 1649977179
transform 1 0 30544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _396_
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _397__37
timestamp 1649977179
transform 1 0 30176 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _397_
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _398__38
timestamp 1649977179
transform 1 0 30820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _398_
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _399__39
timestamp 1649977179
transform 1 0 30820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _399_
timestamp 1649977179
transform 1 0 31832 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _400__40
timestamp 1649977179
transform 1 0 31464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _400_
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _401__41
timestamp 1649977179
transform 1 0 32108 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _401_
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _402__42
timestamp 1649977179
transform 1 0 33764 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _402_
timestamp 1649977179
transform 1 0 34408 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _403__43
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _403_
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _404__44
timestamp 1649977179
transform 1 0 34684 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _404_
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _405__45
timestamp 1649977179
transform 1 0 35972 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _405_
timestamp 1649977179
transform 1 0 34684 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _406__46
timestamp 1649977179
transform 1 0 35972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _406_
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _407__47
timestamp 1649977179
transform 1 0 36156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _407_
timestamp 1649977179
transform 1 0 36984 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _408__48
timestamp 1649977179
transform 1 0 36800 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _408_
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _409__49
timestamp 1649977179
transform 1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _409_
timestamp 1649977179
transform 1 0 37352 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _410__50
timestamp 1649977179
transform 1 0 38180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _410_
timestamp 1649977179
transform 1 0 39560 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _411__51
timestamp 1649977179
transform 1 0 39192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _411_
timestamp 1649977179
transform 1 0 39836 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _412__52
timestamp 1649977179
transform 1 0 39836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _412_
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _413__53
timestamp 1649977179
transform 1 0 40020 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _413_
timestamp 1649977179
transform 1 0 40020 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _414__54
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _414_
timestamp 1649977179
transform 1 0 42412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _415__55
timestamp 1649977179
transform 1 0 41400 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _415_
timestamp 1649977179
transform 1 0 42136 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _416__56
timestamp 1649977179
transform 1 0 43332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _416_
timestamp 1649977179
transform 1 0 42412 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _417__57
timestamp 1649977179
transform 1 0 43056 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _417_
timestamp 1649977179
transform 1 0 42596 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _418__58
timestamp 1649977179
transform 1 0 47564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _418_
timestamp 1649977179
transform 1 0 44712 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _419__59
timestamp 1649977179
transform 1 0 47288 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _419_
timestamp 1649977179
transform 1 0 44988 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _420_
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _420__60
timestamp 1649977179
transform 1 0 47564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _421__61
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _421_
timestamp 1649977179
transform 1 0 44988 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _422__62
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _422_
timestamp 1649977179
transform 1 0 45816 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _423__63
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _423_
timestamp 1649977179
transform 1 0 46276 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _424__64
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _424_
timestamp 1649977179
transform 1 0 45172 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _425__65
timestamp 1649977179
transform 1 0 46184 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _425_
timestamp 1649977179
transform 1 0 45172 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _426__66
timestamp 1649977179
transform 1 0 46920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _426_
timestamp 1649977179
transform 1 0 46276 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _427__67
timestamp 1649977179
transform 1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _427_
timestamp 1649977179
transform 1 0 1564 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _428__68
timestamp 1649977179
transform 1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _428_
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _429__69
timestamp 1649977179
transform 1 0 2392 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _429_
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _430__70
timestamp 1649977179
transform 1 0 3128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _430_
timestamp 1649977179
transform 1 0 1656 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _431__71
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _431_
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _432__72
timestamp 1649977179
transform 1 0 1472 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _432_
timestamp 1649977179
transform 1 0 3956 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _433__73
timestamp 1649977179
transform 1 0 3220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _433_
timestamp 1649977179
transform 1 0 3956 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _434__74
timestamp 1649977179
transform 1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _434_
timestamp 1649977179
transform 1 0 3956 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _435_
timestamp 1649977179
transform 1 0 4232 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _436_
timestamp 1649977179
transform 1 0 6256 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _437_
timestamp 1649977179
transform 1 0 6808 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _438_
timestamp 1649977179
transform 1 0 6532 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _439_
timestamp 1649977179
transform 1 0 6532 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _440_
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _441_
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _442_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _443_
timestamp 1649977179
transform 1 0 6808 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1649977179
transform 1 0 1840 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1649977179
transform 1 0 21804 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1649977179
transform 1 0 25024 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1649977179
transform 1 0 28336 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1649977179
transform 1 0 32108 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1649977179
transform 1 0 34960 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1649977179
transform 1 0 38272 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 42780 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 1649977179
transform 1 0 45356 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 47656 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input11
timestamp 1649977179
transform 1 0 5152 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  repeater12
timestamp 1649977179
transform 1 0 4508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater13
timestamp 1649977179
transform 1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater14
timestamp 1649977179
transform 1 0 10304 0 1 7616
box -38 -48 314 592
<< labels >>
flabel metal2 s 1738 49200 1850 50000 0 FreeSans 448 90 0 0 active
port 0 nsew signal input
flabel metal2 s 21610 49200 21722 50000 0 FreeSans 448 90 0 0 chip_pin_output_bit[0]
port 1 nsew signal input
flabel metal2 s 24922 49200 25034 50000 0 FreeSans 448 90 0 0 chip_pin_output_bit[1]
port 2 nsew signal input
flabel metal2 s 28234 49200 28346 50000 0 FreeSans 448 90 0 0 chip_pin_output_bit[2]
port 3 nsew signal input
flabel metal2 s 31546 49200 31658 50000 0 FreeSans 448 90 0 0 chip_pin_output_bit[3]
port 4 nsew signal input
flabel metal2 s 34858 49200 34970 50000 0 FreeSans 448 90 0 0 chip_pin_output_bit[4]
port 5 nsew signal input
flabel metal2 s 38170 49200 38282 50000 0 FreeSans 448 90 0 0 chip_pin_output_bit[5]
port 6 nsew signal input
flabel metal2 s 41482 49200 41594 50000 0 FreeSans 448 90 0 0 chip_pin_output_bit[6]
port 7 nsew signal input
flabel metal2 s 44794 49200 44906 50000 0 FreeSans 448 90 0 0 chip_pin_output_bit[7]
port 8 nsew signal input
flabel metal2 s 48106 49200 48218 50000 0 FreeSans 448 90 0 0 clk_blip
port 9 nsew signal input
flabel metal3 s 0 3756 800 3996 0 FreeSans 960 0 0 0 io_in[0]
port 10 nsew signal input
flabel metal2 s 11674 49200 11786 50000 0 FreeSans 448 90 0 0 io_in[10]
port 11 nsew signal input
flabel metal2 s 14986 49200 15098 50000 0 FreeSans 448 90 0 0 io_in[11]
port 12 nsew signal input
flabel metal2 s 18298 49200 18410 50000 0 FreeSans 448 90 0 0 io_in[12]
port 13 nsew signal input
flabel metal3 s 0 14636 800 14876 0 FreeSans 960 0 0 0 io_in[13]
port 14 nsew signal input
flabel metal3 s 0 15996 800 16236 0 FreeSans 960 0 0 0 io_in[14]
port 15 nsew signal input
flabel metal3 s 0 17356 800 17596 0 FreeSans 960 0 0 0 io_in[15]
port 16 nsew signal input
flabel metal3 s 0 18716 800 18956 0 FreeSans 960 0 0 0 io_in[16]
port 17 nsew signal input
flabel metal3 s 0 20076 800 20316 0 FreeSans 960 0 0 0 io_in[17]
port 18 nsew signal input
flabel metal3 s 0 21436 800 21676 0 FreeSans 960 0 0 0 io_in[18]
port 19 nsew signal input
flabel metal3 s 0 22796 800 23036 0 FreeSans 960 0 0 0 io_in[19]
port 20 nsew signal input
flabel metal3 s 0 5116 800 5356 0 FreeSans 960 0 0 0 io_in[1]
port 21 nsew signal input
flabel metal3 s 0 24156 800 24396 0 FreeSans 960 0 0 0 io_in[20]
port 22 nsew signal input
flabel metal3 s 0 25516 800 25756 0 FreeSans 960 0 0 0 io_in[21]
port 23 nsew signal input
flabel metal3 s 0 26876 800 27116 0 FreeSans 960 0 0 0 io_in[22]
port 24 nsew signal input
flabel metal3 s 0 28236 800 28476 0 FreeSans 960 0 0 0 io_in[23]
port 25 nsew signal input
flabel metal3 s 0 29596 800 29836 0 FreeSans 960 0 0 0 io_in[24]
port 26 nsew signal input
flabel metal3 s 0 30956 800 31196 0 FreeSans 960 0 0 0 io_in[25]
port 27 nsew signal input
flabel metal3 s 0 32316 800 32556 0 FreeSans 960 0 0 0 io_in[26]
port 28 nsew signal input
flabel metal3 s 0 33676 800 33916 0 FreeSans 960 0 0 0 io_in[27]
port 29 nsew signal input
flabel metal3 s 0 35036 800 35276 0 FreeSans 960 0 0 0 io_in[28]
port 30 nsew signal input
flabel metal3 s 0 36396 800 36636 0 FreeSans 960 0 0 0 io_in[29]
port 31 nsew signal input
flabel metal3 s 0 6476 800 6716 0 FreeSans 960 0 0 0 io_in[2]
port 32 nsew signal input
flabel metal3 s 0 37756 800 37996 0 FreeSans 960 0 0 0 io_in[30]
port 33 nsew signal input
flabel metal3 s 0 39116 800 39356 0 FreeSans 960 0 0 0 io_in[31]
port 34 nsew signal input
flabel metal3 s 0 40476 800 40716 0 FreeSans 960 0 0 0 io_in[32]
port 35 nsew signal input
flabel metal3 s 0 41836 800 42076 0 FreeSans 960 0 0 0 io_in[33]
port 36 nsew signal input
flabel metal3 s 0 43196 800 43436 0 FreeSans 960 0 0 0 io_in[34]
port 37 nsew signal input
flabel metal3 s 0 44556 800 44796 0 FreeSans 960 0 0 0 io_in[35]
port 38 nsew signal input
flabel metal3 s 0 45916 800 46156 0 FreeSans 960 0 0 0 io_in[36]
port 39 nsew signal input
flabel metal3 s 0 47276 800 47516 0 FreeSans 960 0 0 0 io_in[37]
port 40 nsew signal input
flabel metal3 s 0 7836 800 8076 0 FreeSans 960 0 0 0 io_in[3]
port 41 nsew signal input
flabel metal3 s 0 9196 800 9436 0 FreeSans 960 0 0 0 io_in[4]
port 42 nsew signal input
flabel metal3 s 0 10556 800 10796 0 FreeSans 960 0 0 0 io_in[5]
port 43 nsew signal input
flabel metal3 s 0 11916 800 12156 0 FreeSans 960 0 0 0 io_in[6]
port 44 nsew signal input
flabel metal3 s 0 13276 800 13516 0 FreeSans 960 0 0 0 io_in[7]
port 45 nsew signal input
flabel metal2 s 5050 49200 5162 50000 0 FreeSans 448 90 0 0 io_in[8]
port 46 nsew signal input
flabel metal2 s 8362 49200 8474 50000 0 FreeSans 448 90 0 0 io_in[9]
port 47 nsew signal input
flabel metal2 s 25198 0 25310 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 48 nsew signal tristate
flabel metal2 s 31638 0 31750 800 0 FreeSans 448 90 0 0 io_oeb[10]
port 49 nsew signal tristate
flabel metal2 s 32282 0 32394 800 0 FreeSans 448 90 0 0 io_oeb[11]
port 50 nsew signal tristate
flabel metal2 s 32926 0 33038 800 0 FreeSans 448 90 0 0 io_oeb[12]
port 51 nsew signal tristate
flabel metal2 s 33570 0 33682 800 0 FreeSans 448 90 0 0 io_oeb[13]
port 52 nsew signal tristate
flabel metal2 s 34214 0 34326 800 0 FreeSans 448 90 0 0 io_oeb[14]
port 53 nsew signal tristate
flabel metal2 s 34858 0 34970 800 0 FreeSans 448 90 0 0 io_oeb[15]
port 54 nsew signal tristate
flabel metal2 s 35502 0 35614 800 0 FreeSans 448 90 0 0 io_oeb[16]
port 55 nsew signal tristate
flabel metal2 s 36146 0 36258 800 0 FreeSans 448 90 0 0 io_oeb[17]
port 56 nsew signal tristate
flabel metal2 s 36790 0 36902 800 0 FreeSans 448 90 0 0 io_oeb[18]
port 57 nsew signal tristate
flabel metal2 s 37434 0 37546 800 0 FreeSans 448 90 0 0 io_oeb[19]
port 58 nsew signal tristate
flabel metal2 s 25842 0 25954 800 0 FreeSans 448 90 0 0 io_oeb[1]
port 59 nsew signal tristate
flabel metal2 s 38078 0 38190 800 0 FreeSans 448 90 0 0 io_oeb[20]
port 60 nsew signal tristate
flabel metal2 s 38722 0 38834 800 0 FreeSans 448 90 0 0 io_oeb[21]
port 61 nsew signal tristate
flabel metal2 s 39366 0 39478 800 0 FreeSans 448 90 0 0 io_oeb[22]
port 62 nsew signal tristate
flabel metal2 s 40010 0 40122 800 0 FreeSans 448 90 0 0 io_oeb[23]
port 63 nsew signal tristate
flabel metal2 s 40654 0 40766 800 0 FreeSans 448 90 0 0 io_oeb[24]
port 64 nsew signal tristate
flabel metal2 s 41298 0 41410 800 0 FreeSans 448 90 0 0 io_oeb[25]
port 65 nsew signal tristate
flabel metal2 s 41942 0 42054 800 0 FreeSans 448 90 0 0 io_oeb[26]
port 66 nsew signal tristate
flabel metal2 s 42586 0 42698 800 0 FreeSans 448 90 0 0 io_oeb[27]
port 67 nsew signal tristate
flabel metal2 s 43230 0 43342 800 0 FreeSans 448 90 0 0 io_oeb[28]
port 68 nsew signal tristate
flabel metal2 s 43874 0 43986 800 0 FreeSans 448 90 0 0 io_oeb[29]
port 69 nsew signal tristate
flabel metal2 s 26486 0 26598 800 0 FreeSans 448 90 0 0 io_oeb[2]
port 70 nsew signal tristate
flabel metal2 s 44518 0 44630 800 0 FreeSans 448 90 0 0 io_oeb[30]
port 71 nsew signal tristate
flabel metal2 s 45162 0 45274 800 0 FreeSans 448 90 0 0 io_oeb[31]
port 72 nsew signal tristate
flabel metal2 s 45806 0 45918 800 0 FreeSans 448 90 0 0 io_oeb[32]
port 73 nsew signal tristate
flabel metal2 s 46450 0 46562 800 0 FreeSans 448 90 0 0 io_oeb[33]
port 74 nsew signal tristate
flabel metal2 s 47094 0 47206 800 0 FreeSans 448 90 0 0 io_oeb[34]
port 75 nsew signal tristate
flabel metal2 s 47738 0 47850 800 0 FreeSans 448 90 0 0 io_oeb[35]
port 76 nsew signal tristate
flabel metal2 s 48382 0 48494 800 0 FreeSans 448 90 0 0 io_oeb[36]
port 77 nsew signal tristate
flabel metal2 s 49026 0 49138 800 0 FreeSans 448 90 0 0 io_oeb[37]
port 78 nsew signal tristate
flabel metal2 s 27130 0 27242 800 0 FreeSans 448 90 0 0 io_oeb[3]
port 79 nsew signal tristate
flabel metal2 s 27774 0 27886 800 0 FreeSans 448 90 0 0 io_oeb[4]
port 80 nsew signal tristate
flabel metal2 s 28418 0 28530 800 0 FreeSans 448 90 0 0 io_oeb[5]
port 81 nsew signal tristate
flabel metal2 s 29062 0 29174 800 0 FreeSans 448 90 0 0 io_oeb[6]
port 82 nsew signal tristate
flabel metal2 s 29706 0 29818 800 0 FreeSans 448 90 0 0 io_oeb[7]
port 83 nsew signal tristate
flabel metal2 s 30350 0 30462 800 0 FreeSans 448 90 0 0 io_oeb[8]
port 84 nsew signal tristate
flabel metal2 s 30994 0 31106 800 0 FreeSans 448 90 0 0 io_oeb[9]
port 85 nsew signal tristate
flabel metal2 s 726 0 838 800 0 FreeSans 448 90 0 0 io_out[0]
port 86 nsew signal tristate
flabel metal2 s 7166 0 7278 800 0 FreeSans 448 90 0 0 io_out[10]
port 87 nsew signal tristate
flabel metal2 s 7810 0 7922 800 0 FreeSans 448 90 0 0 io_out[11]
port 88 nsew signal tristate
flabel metal2 s 8454 0 8566 800 0 FreeSans 448 90 0 0 io_out[12]
port 89 nsew signal tristate
flabel metal2 s 9098 0 9210 800 0 FreeSans 448 90 0 0 io_out[13]
port 90 nsew signal tristate
flabel metal2 s 9742 0 9854 800 0 FreeSans 448 90 0 0 io_out[14]
port 91 nsew signal tristate
flabel metal2 s 10386 0 10498 800 0 FreeSans 448 90 0 0 io_out[15]
port 92 nsew signal tristate
flabel metal2 s 11030 0 11142 800 0 FreeSans 448 90 0 0 io_out[16]
port 93 nsew signal tristate
flabel metal2 s 11674 0 11786 800 0 FreeSans 448 90 0 0 io_out[17]
port 94 nsew signal tristate
flabel metal2 s 12318 0 12430 800 0 FreeSans 448 90 0 0 io_out[18]
port 95 nsew signal tristate
flabel metal2 s 12962 0 13074 800 0 FreeSans 448 90 0 0 io_out[19]
port 96 nsew signal tristate
flabel metal2 s 1370 0 1482 800 0 FreeSans 448 90 0 0 io_out[1]
port 97 nsew signal tristate
flabel metal2 s 13606 0 13718 800 0 FreeSans 448 90 0 0 io_out[20]
port 98 nsew signal tristate
flabel metal2 s 14250 0 14362 800 0 FreeSans 448 90 0 0 io_out[21]
port 99 nsew signal tristate
flabel metal2 s 14894 0 15006 800 0 FreeSans 448 90 0 0 io_out[22]
port 100 nsew signal tristate
flabel metal2 s 15538 0 15650 800 0 FreeSans 448 90 0 0 io_out[23]
port 101 nsew signal tristate
flabel metal2 s 16182 0 16294 800 0 FreeSans 448 90 0 0 io_out[24]
port 102 nsew signal tristate
flabel metal2 s 16826 0 16938 800 0 FreeSans 448 90 0 0 io_out[25]
port 103 nsew signal tristate
flabel metal2 s 17470 0 17582 800 0 FreeSans 448 90 0 0 io_out[26]
port 104 nsew signal tristate
flabel metal2 s 18114 0 18226 800 0 FreeSans 448 90 0 0 io_out[27]
port 105 nsew signal tristate
flabel metal2 s 18758 0 18870 800 0 FreeSans 448 90 0 0 io_out[28]
port 106 nsew signal tristate
flabel metal2 s 19402 0 19514 800 0 FreeSans 448 90 0 0 io_out[29]
port 107 nsew signal tristate
flabel metal2 s 2014 0 2126 800 0 FreeSans 448 90 0 0 io_out[2]
port 108 nsew signal tristate
flabel metal2 s 20046 0 20158 800 0 FreeSans 448 90 0 0 io_out[30]
port 109 nsew signal tristate
flabel metal2 s 20690 0 20802 800 0 FreeSans 448 90 0 0 io_out[31]
port 110 nsew signal tristate
flabel metal2 s 21334 0 21446 800 0 FreeSans 448 90 0 0 io_out[32]
port 111 nsew signal tristate
flabel metal2 s 21978 0 22090 800 0 FreeSans 448 90 0 0 io_out[33]
port 112 nsew signal tristate
flabel metal2 s 22622 0 22734 800 0 FreeSans 448 90 0 0 io_out[34]
port 113 nsew signal tristate
flabel metal2 s 23266 0 23378 800 0 FreeSans 448 90 0 0 io_out[35]
port 114 nsew signal tristate
flabel metal2 s 23910 0 24022 800 0 FreeSans 448 90 0 0 io_out[36]
port 115 nsew signal tristate
flabel metal2 s 24554 0 24666 800 0 FreeSans 448 90 0 0 io_out[37]
port 116 nsew signal tristate
flabel metal2 s 2658 0 2770 800 0 FreeSans 448 90 0 0 io_out[3]
port 117 nsew signal tristate
flabel metal2 s 3302 0 3414 800 0 FreeSans 448 90 0 0 io_out[4]
port 118 nsew signal tristate
flabel metal2 s 3946 0 4058 800 0 FreeSans 448 90 0 0 io_out[5]
port 119 nsew signal tristate
flabel metal2 s 4590 0 4702 800 0 FreeSans 448 90 0 0 io_out[6]
port 120 nsew signal tristate
flabel metal2 s 5234 0 5346 800 0 FreeSans 448 90 0 0 io_out[7]
port 121 nsew signal tristate
flabel metal2 s 5878 0 5990 800 0 FreeSans 448 90 0 0 io_out[8]
port 122 nsew signal tristate
flabel metal2 s 6522 0 6634 800 0 FreeSans 448 90 0 0 io_out[9]
port 123 nsew signal tristate
flabel metal4 s 4208 2128 4528 47376 0 FreeSans 1920 90 0 0 vccd1
port 124 nsew power bidirectional
flabel metal4 s 34928 2128 35248 47376 0 FreeSans 1920 90 0 0 vccd1
port 124 nsew power bidirectional
flabel metal4 s 19568 2128 19888 47376 0 FreeSans 1920 90 0 0 vssd1
port 125 nsew ground bidirectional
flabel metal3 s 0 2396 800 2636 0 FreeSans 960 0 0 0 wb_clk_i
port 126 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
